----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 07/29/2020 03:02:34 PM
-- Design Name: 
-- Module Name: input_ram - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity input_ram is
Port ( clk : in  STD_LOGIC;
           cs : in  STD_LOGIC;
         --  we : in  STD_LOGIC;

           address : in integer;-- range 0 to 65535;--STD_LOGIC_VECTOR(2 downto 0);
           data_out : out  integer range 0 to 255);--STD_LOGIC_VECTOR (63 downto 0));
end input_ram;

architecture Behavioral of input_ram is

type mem_array is array(65535 downto 0)  of integer range 0 to 255;--std_logic_vector(63 downto 0);

--constant memory:MEM_array:=(150, 144, 155, 157, 105, 164, 173, 173, 171, 173, 177, 181, 178, 183, 178, 180, 184, 186, 190, 183, 185, 185, 184, 188, 188, 185, 183, 190, 187, 187, 188, 186, 190, 189, 190, 190, 190, 192, 193, 193, 193, 192, 191, 194, 197, 195, 198, 196, 194, 193, 193, 196, 194, 199, 198, 200, 198, 198, 195, 195, 196, 200, 200, 198, 199, 199, 200, 197, 198, 199, 203, 198, 202, 200, 200, 200, 200, 201, 201, 200, 202, 199, 200, 201, 203, 199, 204, 201, 202, 205, 204, 204, 199, 202, 201, 202, 200, 203, 201, 204, 205, 203, 201, 204, 205, 208, 207, 208, 207, 206, 210, 208, 205, 204, 204, 207, 207, 208, 203, 207, 205, 206, 204, 203, 200, 201, 205, 203, 205, 205, 207, 208, 203, 208, 210, 205, 205, 205, 204, 208, 213, 209, 207, 209, 210, 207, 206, 203, 204, 207, 207, 208, 204, 206, 207, 208, 205, 206, 207, 208, 207, 208, 209, 206, 207, 208, 205, 210, 204, 202, 206, 201, 205, 207, 205, 204, 203, 204, 206, 202, 202, 199, 203, 201, 202, 200, 203, 202, 203, 203, 203, 201, 202, 203, 204, 203, 199, 201, 200, 199, 200, 201, 201, 198, 202, 197, 202, 204, 198, 204, 214, 204, 198, 199, 200, 201, 201, 199, 195, 198, 198, 200, 198, 197, 192, 198, 199, 199, 193, 200, 200, 197, 195, 196, 194, 195, 197, 192, 195, 195, 195, 195, 196, 192, 194, 195, 193, 191, 190, 194, 193, 190, 186, 189, 188, 161, 189, 183, 185, 184, 112, 185, 182, 184, 185, 187, 184, 192, 188, 192, 184, 188, 188, 188, 192, 193, 194, 192, 193, 190, 195, 189, 190, 192, 192, 192, 193, 191, 195, 197, 195, 196, 194, 195, 196, 197, 191, 194, 196, 196, 197, 196, 192, 198, 194, 192, 196, 195, 197, 199, 197, 200, 197, 199, 197, 197, 197, 199, 201, 196, 201, 201, 204, 202, 200, 201, 205, 197, 199, 205, 203, 200, 199, 204, 205, 199, 205, 203, 204, 203, 202, 201, 202, 203, 203, 206, 205, 203, 203, 203, 200, 207, 205, 205, 206, 207, 204, 206, 202, 206, 209, 209, 212, 209, 209, 208, 212, 213, 208, 204, 205, 208, 207, 206, 208, 207, 209, 208, 211, 209, 202, 204, 206, 205, 209, 208, 206, 206, 208, 209, 209, 207, 206, 208, 208, 211, 214, 212, 210, 209, 208, 209, 206, 208, 205, 206, 208, 209, 208, 209, 207, 208, 211, 211, 208, 207, 209, 207, 206, 208, 204, 207, 209, 210, 206, 207, 205, 208, 206, 210, 207, 203, 204, 207, 205, 204, 208, 204, 204, 206, 204, 204, 203, 206, 204, 205, 203, 198, 202, 207, 203, 205, 200, 200, 198, 200, 204, 200, 200, 197, 200, 197, 200, 198, 197, 198, 199, 201, 202, 204, 202, 203, 202, 198, 199, 198, 197, 200, 199, 197, 194, 197, 199, 200, 200, 196, 195, 201, 197, 197, 193, 191, 195, 192, 196, 198, 198, 198, 197, 200, 199, 193, 194, 191, 192, 192, 192, 190, 188, 185, 185, 121, 191, 184, 183, 189, 115, 183, 184, 185, 190, 188, 185, 188, 186, 190, 187, 190, 190, 194, 191, 189, 194, 193, 191, 191, 192, 193, 189, 190, 193, 196, 193, 192, 194, 198, 190, 191, 196, 194, 195, 198, 193, 196, 195, 197, 197, 196, 195, 199, 194, 190, 195, 196, 197, 198, 199, 199, 200, 200, 194, 198, 197, 197, 199, 202, 198, 204, 204, 200, 202, 204, 203, 202, 201, 206, 200, 204, 202, 205, 204, 204, 205, 202, 202, 207, 202, 206, 200, 204, 203, 212, 207, 205, 204, 203, 206, 206, 209, 207, 207, 210, 208, 205, 205, 205, 209, 207, 210, 209, 208, 210, 209, 212, 206, 208, 205, 208, 208, 208, 208, 206, 205, 208, 207, 208, 207, 204, 206, 208, 206, 210, 209, 209, 209, 212, 209, 207, 206, 206, 208, 211, 213, 212, 208, 209, 209, 207, 208, 206, 207, 205, 208, 209, 207, 207, 210, 213, 207, 209, 208, 207, 208, 210, 210, 207, 205, 208, 208, 208, 208, 206, 209, 204, 204, 207, 206, 209, 203, 207, 201, 201, 207, 205, 205, 205, 206, 205, 201, 205, 204, 205, 203, 198, 204, 206, 204, 206, 201, 202, 204, 204, 204, 203, 199, 196, 201, 199, 204, 200, 201, 199, 200, 204, 202, 203, 199, 204, 203, 202, 200, 202, 203, 199, 203, 203, 199, 196, 198, 200, 200, 201, 197, 202, 197, 194, 199, 196, 195, 194, 200, 200, 200, 198, 197, 199, 198, 193, 195, 192, 194, 192, 194, 190, 188, 189, 183, 113, 189, 186, 183, 189, 113, 182, 185, 187, 187, 188, 184, 185, 190, 188, 189, 190, 192, 191, 193, 196, 195, 196, 194, 192, 191, 194, 190, 191, 198, 189, 193, 191, 192, 196, 193, 191, 193, 192, 193, 199, 197, 195, 197, 198, 201, 199, 200, 196, 199, 196, 198, 198, 201, 198, 198, 199, 200, 202, 198, 203, 198, 200, 201, 203, 202, 205, 201, 204, 201, 199, 199, 199, 200, 201, 203, 200, 201, 206, 205, 205, 203, 205, 208, 204, 207, 206, 200, 205, 204, 208, 205, 201, 204, 205, 204, 205, 208, 209, 209, 209, 209, 204, 205, 206, 207, 211, 210, 207, 208, 205, 209, 210, 209, 207, 206, 209, 209, 207, 211, 207, 206, 206, 208, 208, 206, 206, 210, 209, 208, 210, 209, 208, 209, 209, 208, 206, 206, 211, 212, 212, 214, 211, 208, 209, 209, 208, 207, 202, 207, 208, 210, 208, 208, 210, 208, 210, 211, 208, 205, 205, 210, 210, 212, 209, 209, 205, 208, 209, 205, 206, 207, 202, 207, 205, 206, 205, 204, 208, 202, 206, 207, 206, 207, 205, 204, 201, 205, 205, 205, 206, 202, 198, 203, 203, 206, 208, 201, 203, 204, 205, 203, 202, 200, 199, 202, 202, 200, 198, 204, 199, 200, 204, 203, 205, 201, 200, 203, 203, 204, 204, 203, 203, 202, 202, 200, 199, 198, 201, 199, 198, 198, 202, 199, 197, 195, 197, 198, 194, 197, 196, 199, 194, 195, 199, 195, 194, 195, 193, 196, 195, 189, 194, 184, 185, 182, 115, 186, 182, 180, 189, 120, 187, 189, 187, 188, 182, 185, 184, 184, 185, 186, 191, 188, 192, 196, 195, 195, 198, 193, 189, 191, 192, 193, 190, 193, 192, 194, 192, 192, 195, 191, 194, 190, 191, 194, 198, 198, 195, 198, 197, 203, 201, 199, 195, 195, 198, 198, 198, 201, 200, 199, 200, 198, 196, 197, 201, 198, 201, 200, 198, 202, 203, 201, 201, 204, 199, 201, 201, 201, 202, 206, 206, 201, 205, 205, 207, 205, 204, 206, 204, 204, 203, 200, 200, 203, 205, 204, 203, 203, 206, 207, 206, 208, 207, 207, 207, 208, 204, 203, 207, 208, 209, 211, 210, 206, 209, 210, 211, 208, 207, 206, 211, 211, 205, 210, 206, 207, 212, 206, 208, 208, 204, 206, 205, 207, 210, 209, 208, 207, 208, 207, 209, 212, 211, 212, 212, 214, 210, 210, 213, 210, 210, 208, 207, 208, 209, 211, 209, 210, 213, 209, 210, 209, 212, 207, 205, 209, 212, 208, 209, 210, 207, 208, 209, 207, 209, 208, 205, 207, 208, 205, 208, 204, 206, 206, 208, 208, 207, 206, 204, 210, 203, 206, 204, 203, 204, 203, 200, 203, 207, 204, 205, 204, 205, 205, 203, 204, 206, 200, 200, 202, 202, 204, 201, 202, 203, 200, 206, 203, 206, 204, 202, 203, 204, 205, 200, 199, 200, 202, 204, 199, 203, 197, 200, 198, 197, 205, 199, 203, 196, 199, 197, 197, 198, 197, 198, 202, 195, 197, 196, 193, 197, 195, 195, 193, 198, 196, 193, 190, 188, 186, 131, 187, 185, 187, 192, 107, 184, 193, 192, 185, 188, 185, 187, 185, 188, 188, 188, 189, 193, 194, 195, 195, 193, 193, 191, 195, 193, 191, 192, 194, 192, 193, 192, 192, 194, 194, 195, 195, 192, 197, 196, 201, 197, 194, 198, 200, 201, 199, 198, 198, 198, 199, 198, 199, 200, 194, 199, 194, 197, 200, 202, 203, 201, 201, 202, 203, 202, 201, 202, 202, 200, 200, 202, 203, 206, 205, 203, 204, 208, 210, 208, 204, 202, 204, 200, 202, 200, 200, 199, 202, 204, 205, 206, 205, 205, 206, 207, 209, 208, 207, 209, 206, 207, 205, 207, 209, 208, 208, 209, 209, 210, 208, 209, 211, 208, 208, 208, 211, 208, 204, 206, 204, 207, 207, 204, 205, 208, 210, 211, 209, 208, 207, 208, 207, 209, 210, 210, 214, 212, 211, 209, 211, 208, 208, 210, 207, 211, 207, 209, 208, 206, 216, 215, 212, 211, 210, 213, 207, 214, 206, 208, 209, 211, 210, 213, 211, 210, 211, 206, 210, 211, 206, 204, 210, 206, 203, 205, 205, 206, 205, 208, 206, 204, 208, 207, 206, 206, 204, 204, 203, 206, 203, 201, 205, 204, 206, 208, 204, 202, 204, 203, 202, 206, 200, 203, 204, 201, 203, 203, 204, 202, 202, 200, 202, 206, 200, 203, 202, 202, 202, 202, 199, 202, 202, 200, 203, 202, 203, 205, 197, 199, 202, 198, 201, 200, 200, 195, 197, 197, 197, 200, 197, 197, 195, 196, 193, 196, 198, 200, 198, 198, 198, 193, 195, 187, 181, 119, 190, 188, 186, 190, 115, 184, 190, 188, 189, 185, 183, 185, 184, 188, 186, 190, 192, 194, 194, 198, 194, 193, 194, 194, 192, 190, 189, 189, 192, 193, 192, 193, 190, 193, 196, 195, 194, 193, 195, 200, 199, 193, 198, 199, 197, 200, 199, 199, 199, 196, 203, 197, 199, 198, 197, 198, 200, 201, 197, 204, 204, 204, 203, 200, 200, 202, 204, 203, 200, 201, 201, 204, 203, 205, 205, 203, 208, 207, 209, 208, 203, 200, 204, 204, 203, 201, 202, 203, 205, 205, 207, 206, 206, 207, 207, 210, 209, 209, 208, 209, 206, 204, 204, 205, 207, 207, 211, 208, 210, 207, 210, 207, 210, 207, 210, 207, 210, 208, 207, 206, 205, 209, 210, 204, 203, 204, 204, 207, 208, 207, 212, 211, 211, 207, 212, 207, 212, 210, 209, 209, 213, 208, 209, 210, 211, 211, 207, 212, 210, 211, 210, 213, 211, 209, 208, 212, 210, 211, 209, 208, 210, 212, 212, 208, 210, 213, 209, 209, 212, 209, 205, 207, 209, 209, 207, 207, 208, 206, 205, 206, 208, 208, 206, 208, 206, 209, 208, 204, 207, 211, 203, 207, 206, 207, 208, 207, 203, 204, 206, 208, 206, 204, 208, 203, 205, 202, 203, 201, 201, 203, 205, 204, 204, 202, 201, 203, 203, 203, 204, 200, 203, 205, 203, 207, 203, 203, 200, 204, 200, 200, 202, 200, 202, 199, 201, 199, 199, 194, 196, 193, 192, 192, 193, 196, 195, 195, 194, 196, 195, 197, 198, 196, 192, 189, 182, 106, 189, 184, 185, 188, 102, 184, 191, 191, 183, 186, 185, 188, 183, 186, 188, 190, 189, 189, 195, 195, 196, 190, 191, 193, 187, 189, 192, 191, 191, 197, 192, 195, 193, 197, 197, 192, 194, 197, 197, 201, 197, 198, 198, 197, 201, 201, 201, 199, 198, 198, 201, 201, 197, 201, 199, 200, 199, 199, 201, 201, 201, 205, 203, 201, 203, 200, 206, 201, 204, 203, 206, 204, 205, 204, 202, 204, 205, 208, 206, 207, 204, 201, 203, 201, 202, 204, 205, 207, 210, 205, 206, 204, 206, 206, 207, 211, 211, 207, 207, 211, 207, 207, 208, 207, 210, 209, 209, 209, 209, 206, 211, 207, 207, 209, 208, 205, 211, 209, 209, 203, 204, 206, 209, 206, 209, 205, 207, 204, 207, 207, 211, 209, 208, 208, 207, 208, 209, 210, 211, 211, 213, 211, 210, 211, 211, 211, 211, 210, 211, 212, 210, 207, 213, 211, 212, 210, 211, 211, 211, 209, 212, 211, 215, 208, 210, 209, 211, 212, 210, 210, 208, 207, 208, 208, 208, 208, 205, 205, 208, 207, 207, 209, 209, 206, 208, 210, 207, 209, 206, 207, 207, 206, 207, 208, 209, 208, 208, 203, 209, 203, 208, 209, 205, 203, 204, 204, 202, 202, 201, 202, 201, 202, 203, 199, 203, 202, 205, 209, 208, 201, 204, 205, 207, 207, 206, 204, 201, 205, 202, 201, 202, 201, 199, 200, 200, 197, 201, 199, 197, 198, 199, 193, 196, 202, 200, 196, 196, 199, 198, 199, 201, 196, 192, 192, 183, 107, 185, 185, 182, 186, 117, 187, 191, 191, 185, 191, 184, 188, 186, 188, 189, 189, 189, 196, 195, 192, 193, 194, 193, 195, 195, 193, 192, 194, 193, 194, 194, 193, 195, 198, 194, 197, 197, 193, 196, 200, 199, 200, 201, 200, 205, 200, 199, 203, 201, 196, 200, 201, 200, 197, 199, 201, 203, 201, 201, 204, 201, 206, 205, 202, 204, 204, 206, 203, 207, 203, 204, 202, 204, 204, 203, 197, 201, 207, 208, 209, 205, 205, 202, 205, 205, 206, 206, 208, 210, 207, 207, 204, 206, 208, 210, 212, 210, 208, 205, 206, 208, 207, 207, 209, 210, 210, 208, 207, 205, 209, 210, 210, 208, 207, 207, 209, 208, 207, 207, 209, 208, 212, 206, 207, 206, 207, 208, 203, 202, 207, 207, 208, 209, 207, 202, 203, 206, 207, 213, 211, 214, 211, 208, 213, 211, 212, 212, 211, 208, 212, 212, 209, 211, 210, 211, 210, 210, 210, 208, 211, 209, 213, 210, 209, 208, 210, 208, 210, 211, 211, 207, 204, 209, 208, 208, 206, 211, 209, 206, 207, 204, 203, 207, 206, 209, 206, 203, 208, 206, 205, 205, 208, 209, 209, 208, 209, 207, 203, 207, 208, 207, 205, 206, 206, 208, 205, 201, 203, 202, 204, 204, 203, 207, 203, 201, 203, 203, 207, 206, 203, 208, 209, 206, 210, 205, 203, 206, 206, 203, 202, 200, 200, 201, 200, 202, 198, 198, 198, 197, 197, 197, 194, 195, 201, 202, 197, 199, 203, 201, 203, 200, 199, 196, 193, 188, 114, 188, 186, 178, 191, 116, 185, 190, 194, 188, 192, 187, 191, 186, 185, 190, 186, 190, 192, 193, 193, 192, 192, 195, 195, 190, 196, 195, 191, 197, 196, 192, 195, 194, 196, 195, 198, 196, 197, 200, 203, 200, 199, 201, 200, 203, 203, 203, 203, 204, 199, 200, 204, 202, 195, 197, 200, 202, 202, 204, 203, 202, 205, 204, 203, 201, 205, 205, 206, 206, 203, 204, 203, 207, 207, 205, 197, 198, 207, 210, 210, 206, 205, 201, 207, 202, 208, 207, 205, 210, 209, 207, 208, 205, 210, 208, 211, 210, 207, 205, 213, 210, 210, 206, 209, 212, 208, 210, 210, 205, 209, 214, 211, 210, 209, 207, 207, 208, 210, 208, 208, 208, 207, 205, 206, 207, 207, 206, 206, 209, 208, 206, 210, 207, 205, 203, 206, 210, 211, 213, 213, 213, 212, 210, 209, 209, 209, 211, 213, 210, 212, 212, 209, 205, 205, 207, 208, 210, 212, 208, 211, 210, 208, 212, 207, 206, 213, 207, 209, 203, 206, 204, 206, 212, 210, 208, 205, 209, 207, 208, 208, 206, 204, 207, 206, 208, 211, 208, 210, 207, 210, 206, 203, 211, 209, 209, 207, 206, 205, 205, 203, 208, 206, 206, 203, 209, 204, 203, 203, 202, 204, 206, 202, 203, 202, 201, 201, 203, 206, 207, 207, 209, 209, 210, 208, 207, 204, 203, 203, 203, 204, 199, 202, 204, 200, 203, 200, 198, 202, 202, 199, 196, 197, 196, 199, 199, 199, 197, 201, 201, 202, 197, 200, 195, 196, 188, 122, 188, 186, 187, 188, 105, 189, 193, 191, 185, 190, 189, 195, 192, 189, 186, 188, 191, 195, 194, 193, 189, 197, 192, 195, 198, 194, 200, 200, 196, 192, 192, 195, 194, 197, 196, 196, 199, 198, 199, 202, 202, 202, 199, 200, 203, 204, 201, 200, 202, 201, 201, 203, 200, 197, 197, 200, 203, 204, 206, 204, 203, 206, 203, 205, 202, 202, 206, 208, 205, 204, 202, 202, 206, 205, 204, 207, 207, 207, 209, 209, 204, 204, 202, 205, 207, 210, 208, 207, 206, 205, 206, 206, 207, 207, 209, 208, 213, 209, 210, 213, 211, 210, 203, 207, 207, 207, 209, 213, 212, 208, 211, 216, 210, 211, 210, 208, 210, 210, 208, 209, 206, 206, 208, 202, 203, 205, 205, 206, 209, 208, 206, 209, 210, 210, 205, 206, 212, 210, 212, 216, 215, 214, 211, 212, 210, 211, 211, 208, 214, 213, 213, 210, 206, 209, 207, 208, 213, 211, 211, 212, 209, 213, 210, 212, 213, 214, 208, 208, 210, 206, 210, 209, 210, 211, 210, 209, 207, 209, 210, 209, 207, 208, 208, 208, 208, 205, 207, 204, 207, 209, 208, 205, 208, 205, 209, 209, 208, 204, 205, 206, 208, 206, 205, 203, 206, 207, 206, 205, 205, 205, 209, 204, 207, 201, 204, 199, 205, 208, 207, 207, 204, 209, 208, 207, 206, 206, 203, 207, 204, 200, 203, 197, 203, 206, 203, 200, 206, 204, 205, 203, 196, 195, 199, 197, 200, 200, 199, 202, 201, 204, 198, 202, 202, 195, 192, 134, 190, 184, 186, 186, 116, 186, 193, 188, 186, 187, 188, 192, 193, 192, 190, 189, 193, 191, 195, 194, 195, 197, 196, 196, 197, 196, 198, 200, 195, 198, 196, 199, 196, 199, 199, 198, 198, 196, 200, 202, 201, 201, 201, 204, 204, 201, 202, 201, 204, 203, 206, 203, 202, 201, 199, 201, 207, 206, 203, 203, 202, 206, 207, 202, 207, 203, 204, 205, 206, 204, 205, 204, 207, 202, 206, 205, 208, 209, 209, 205, 207, 201, 204, 204, 207, 211, 208, 207, 209, 206, 208, 206, 208, 205, 211, 210, 212, 213, 213, 213, 214, 212, 208, 208, 207, 210, 212, 214, 213, 212, 212, 215, 214, 216, 212, 208, 210, 210, 207, 208, 204, 204, 209, 204, 207, 204, 204, 206, 210, 212, 209, 211, 209, 212, 210, 207, 210, 213, 212, 217, 212, 210, 211, 206, 210, 210, 213, 213, 212, 212, 216, 213, 209, 210, 212, 211, 215, 212, 210, 207, 209, 211, 211, 213, 214, 214, 212, 211, 211, 208, 208, 209, 212, 210, 210, 207, 210, 211, 210, 207, 208, 205, 211, 212, 209, 209, 206, 206, 210, 205, 207, 207, 206, 205, 209, 207, 208, 206, 204, 204, 205, 206, 203, 207, 207, 207, 206, 208, 208, 205, 210, 207, 209, 205, 204, 204, 201, 206, 203, 204, 208, 205, 204, 207, 208, 203, 206, 205, 205, 202, 205, 200, 205, 207, 200, 202, 202, 204, 205, 204, 198, 199, 198, 200, 201, 200, 199, 204, 207, 201, 203, 201, 201, 199, 190, 127, 187, 185, 186, 192, 104, 194, 192, 189, 188, 188, 186, 184, 192, 190, 188, 192, 191, 192, 192, 195, 195, 195, 194, 198, 199, 196, 197, 197, 197, 196, 198, 198, 196, 196, 196, 196, 194, 199, 198, 200, 199, 202, 202, 201, 206, 201, 205, 202, 201, 201, 203, 200, 198, 198, 198, 201, 204, 206, 201, 204, 205, 204, 209, 204, 205, 206, 209, 207, 208, 207, 205, 205, 205, 204, 205, 205, 207, 208, 209, 205, 206, 204, 206, 207, 206, 207, 206, 209, 208, 209, 211, 210, 205, 207, 207, 212, 209, 209, 213, 212, 211, 211, 209, 207, 209, 210, 209, 212, 210, 211, 213, 211, 212, 211, 211, 209, 208, 207, 209, 211, 208, 207, 207, 206, 203, 207, 202, 205, 209, 208, 207, 209, 211, 211, 208, 208, 210, 214, 212, 214, 212, 212, 214, 208, 210, 213, 213, 210, 211, 214, 214, 212, 208, 211, 214, 211, 212, 212, 208, 211, 209, 210, 210, 211, 212, 211, 210, 210, 212, 209, 208, 210, 210, 212, 211, 209, 210, 212, 211, 210, 209, 205, 210, 209, 207, 208, 206, 208, 211, 208, 209, 207, 207, 211, 208, 210, 211, 205, 207, 207, 205, 206, 208, 207, 206, 211, 208, 206, 207, 206, 206, 208, 207, 209, 205, 202, 204, 203, 203, 207, 207, 205, 209, 210, 206, 206, 210, 206, 205, 203, 201, 205, 201, 204, 206, 205, 204, 208, 205, 201, 198, 201, 199, 198, 201, 204, 199, 201, 205, 202, 203, 201, 200, 198, 193, 141, 188, 186, 183, 188, 109, 187, 190, 185, 189, 193, 189, 188, 194, 192, 190, 192, 193, 192, 193, 192, 195, 193, 197, 196, 202, 197, 198, 196, 194, 199, 199, 199, 197, 199, 192, 200, 197, 200, 199, 197, 199, 204, 201, 203, 205, 204, 202, 204, 200, 205, 203, 204, 197, 197, 200, 203, 205, 203, 203, 205, 202, 205, 209, 206, 205, 206, 208, 205, 206, 205, 204, 204, 206, 205, 203, 204, 204, 205, 207, 208, 206, 208, 207, 209, 207, 208, 208, 208, 211, 210, 211, 210, 207, 209, 208, 210, 208, 209, 211, 213, 213, 209, 209, 211, 211, 208, 208, 211, 212, 210, 213, 216, 215, 212, 212, 212, 212, 210, 207, 210, 209, 209, 207, 209, 205, 208, 204, 201, 207, 207, 211, 210, 206, 213, 207, 207, 213, 211, 214, 213, 210, 209, 212, 210, 213, 211, 211, 212, 212, 213, 211, 209, 211, 213, 211, 213, 214, 215, 211, 212, 214, 211, 212, 210, 212, 209, 211, 208, 210, 210, 207, 211, 212, 211, 211, 213, 212, 212, 211, 206, 208, 206, 212, 209, 210, 208, 208, 211, 208, 210, 211, 207, 207, 208, 207, 209, 209, 210, 209, 206, 205, 208, 208, 208, 208, 206, 209, 207, 207, 207, 205, 206, 205, 209, 205, 206, 203, 209, 207, 207, 208, 210, 208, 209, 208, 207, 208, 203, 207, 200, 204, 206, 202, 206, 210, 206, 205, 206, 204, 202, 201, 199, 198, 198, 202, 201, 195, 201, 202, 204, 204, 207, 201, 195, 191, 144, 192, 187, 183, 187, 107, 190, 192, 190, 188, 189, 187, 191, 192, 193, 196, 188, 195, 196, 197, 194, 191, 198, 199, 195, 198, 196, 198, 197, 196, 196, 198, 196, 198, 198, 196, 198, 197, 197, 197, 198, 201, 201, 205, 205, 205, 205, 204, 204, 203, 201, 203, 204, 201, 202, 207, 204, 206, 206, 203, 202, 204, 205, 204, 206, 204, 205, 204, 205, 205, 205, 205, 204, 205, 206, 204, 206, 206, 206, 209, 211, 207, 209, 208, 208, 210, 209, 206, 208, 210, 213, 210, 211, 212, 213, 209, 210, 210, 210, 209, 212, 212, 214, 209, 211, 213, 214, 211, 213, 212, 213, 215, 214, 215, 213, 213, 213, 210, 210, 207, 207, 213, 211, 208, 213, 209, 207, 204, 203, 207, 206, 208, 209, 209, 209, 213, 208, 212, 212, 212, 211, 212, 209, 207, 211, 211, 210, 213, 213, 212, 213, 211, 212, 215, 211, 210, 212, 216, 213, 212, 212, 214, 214, 212, 212, 212, 212, 211, 207, 210, 209, 208, 209, 211, 211, 209, 210, 211, 214, 209, 211, 208, 205, 210, 211, 212, 206, 208, 210, 209, 213, 210, 208, 206, 209, 207, 209, 211, 208, 213, 208, 206, 210, 208, 206, 209, 203, 207, 208, 207, 208, 208, 208, 209, 207, 206, 210, 208, 207, 209, 206, 207, 206, 210, 210, 209, 205, 206, 204, 205, 204, 203, 207, 206, 208, 208, 207, 207, 206, 206, 204, 201, 201, 203, 199, 205, 199, 201, 202, 203, 204, 206, 205, 200, 196, 188, 142, 191, 189, 184, 189, 98, 186, 187, 188, 194, 189, 191, 191, 194, 193, 194, 197, 195, 194, 196, 195, 197, 197, 202, 200, 199, 198, 196, 197, 199, 198, 198, 203, 199, 197, 198, 202, 198, 199, 195, 194, 201, 204, 203, 203, 208, 203, 200, 202, 203, 207, 205, 206, 202, 200, 202, 204, 205, 205, 203, 204, 203, 205, 202, 202, 206, 207, 207, 206, 209, 207, 203, 203, 205, 207, 207, 209, 202, 205, 207, 211, 207, 209, 208, 209, 210, 209, 208, 210, 213, 214, 210, 212, 208, 213, 212, 212, 209, 211, 211, 211, 212, 215, 213, 211, 214, 213, 214, 212, 214, 215, 215, 217, 217, 215, 217, 214, 211, 209, 211, 209, 212, 210, 207, 211, 211, 210, 208, 205, 207, 209, 212, 210, 210, 213, 212, 212, 212, 213, 215, 215, 213, 212, 207, 213, 212, 211, 209, 213, 214, 214, 217, 217, 213, 211, 211, 217, 213, 216, 213, 213, 214, 212, 216, 213, 212, 208, 210, 207, 204, 210, 207, 207, 211, 215, 212, 209, 212, 216, 209, 212, 209, 209, 210, 211, 209, 204, 209, 212, 210, 214, 212, 206, 207, 210, 208, 211, 209, 208, 209, 209, 207, 207, 207, 207, 211, 206, 209, 204, 209, 210, 209, 207, 207, 209, 209, 208, 205, 208, 204, 210, 207, 210, 213, 211, 209, 205, 205, 206, 202, 205, 204, 207, 207, 210, 206, 203, 205, 206, 206, 206, 203, 202, 200, 203, 206, 204, 204, 200, 200, 202, 204, 201, 199, 194, 191, 140, 195, 188, 187, 187, 110, 189, 190, 192, 190, 190, 185, 189, 193, 191, 192, 190, 193, 197, 201, 194, 196, 196, 200, 198, 197, 198, 196, 194, 195, 197, 198, 203, 199, 204, 200, 203, 199, 201, 199, 201, 202, 202, 200, 201, 191, 204, 202, 202, 204, 204, 206, 207, 205, 203, 205, 205, 205, 205, 204, 203, 205, 207, 203, 203, 205, 206, 209, 202, 204, 208, 204, 206, 209, 208, 211, 210, 206, 207, 206, 207, 211, 208, 208, 210, 212, 211, 211, 212, 210, 214, 212, 213, 211, 210, 213, 213, 212, 209, 214, 211, 214, 213, 212, 213, 214, 214, 213, 213, 214, 214, 213, 217, 217, 218, 215, 213, 208, 208, 209, 208, 209, 210, 209, 211, 211, 207, 209, 206, 208, 210, 210, 208, 210, 214, 215, 213, 216, 216, 219, 215, 215, 214, 212, 211, 213, 211, 214, 215, 214, 213, 217, 216, 215, 214, 211, 216, 216, 218, 216, 215, 211, 212, 215, 214, 211, 213, 209, 207, 210, 210, 208, 210, 210, 211, 208, 213, 207, 215, 206, 211, 211, 212, 212, 213, 212, 205, 209, 210, 209, 211, 211, 209, 208, 203, 210, 208, 209, 209, 209, 210, 211, 212, 210, 209, 212, 209, 210, 212, 205, 208, 210, 208, 209, 208, 207, 206, 205, 204, 205, 209, 204, 214, 212, 213, 210, 210, 210, 209, 208, 209, 205, 211, 210, 209, 209, 206, 207, 205, 204, 205, 205, 201, 201, 203, 205, 204, 206, 205, 203, 203, 206, 203, 200, 198, 193, 143, 196, 190, 190, 189, 106, 185, 194, 191, 193, 189, 184, 187, 191, 197, 192, 193, 194, 196, 198, 197, 197, 197, 199, 197, 196, 199, 196, 199, 197, 203, 198, 202, 199, 206, 204, 202, 199, 200, 198, 198, 201, 202, 202, 201, 200, 205, 204, 205, 208, 203, 208, 204, 205, 202, 208, 206, 206, 206, 203, 205, 206, 209, 208, 205, 205, 203, 209, 205, 208, 208, 208, 209, 212, 210, 213, 210, 208, 208, 208, 207, 211, 206, 208, 210, 212, 214, 209, 212, 212, 211, 210, 211, 210, 211, 213, 210, 211, 213, 215, 215, 213, 212, 213, 214, 213, 214, 214, 212, 214, 213, 214, 216, 217, 216, 214, 214, 211, 208, 209, 209, 209, 210, 212, 211, 212, 210, 211, 209, 209, 210, 211, 209, 210, 212, 214, 215, 214, 212, 216, 213, 216, 213, 210, 214, 211, 213, 213, 214, 214, 215, 216, 218, 216, 212, 212, 209, 217, 214, 214, 212, 214, 215, 212, 212, 213, 211, 211, 208, 209, 213, 210, 211, 214, 208, 209, 212, 212, 213, 213, 210, 209, 210, 210, 211, 209, 208, 204, 204, 209, 211, 207, 207, 210, 208, 212, 213, 208, 212, 209, 207, 209, 209, 210, 210, 210, 212, 211, 209, 207, 207, 208, 208, 208, 207, 207, 207, 204, 207, 204, 205, 207, 212, 210, 214, 210, 210, 212, 212, 209, 208, 209, 208, 210, 209, 211, 209, 207, 204, 206, 205, 208, 203, 203, 204, 206, 209, 205, 206, 204, 204, 207, 203, 200, 196, 191, 139, 195, 189, 191, 190, 106, 189, 192, 190, 190, 189, 193, 196, 194, 195, 190, 194, 196, 201, 198, 195, 196, 196, 196, 198, 198, 195, 198, 197, 195, 199, 200, 202, 200, 204, 203, 201, 200, 202, 199, 202, 203, 202, 202, 205, 207, 207, 208, 211, 207, 207, 207, 205, 207, 204, 206, 208, 206, 205, 205, 206, 208, 207, 206, 209, 208, 211, 213, 211, 212, 208, 210, 210, 212, 211, 213, 208, 210, 209, 210, 211, 209, 211, 211, 212, 211, 211, 211, 212, 212, 213, 205, 212, 211, 212, 211, 212, 213, 213, 213, 215, 213, 210, 212, 215, 214, 213, 214, 214, 213, 212, 214, 216, 215, 216, 211, 213, 212, 209, 212, 209, 212, 210, 216, 214, 213, 213, 210, 210, 211, 211, 206, 212, 212, 213, 217, 216, 214, 216, 219, 217, 213, 214, 214, 216, 212, 214, 216, 213, 215, 219, 218, 217, 216, 209, 212, 212, 215, 214, 216, 215, 214, 217, 214, 214, 211, 212, 211, 211, 214, 212, 212, 211, 213, 210, 213, 211, 210, 211, 215, 214, 211, 209, 211, 209, 210, 205, 206, 206, 210, 210, 214, 209, 209, 207, 210, 211, 208, 208, 210, 210, 210, 212, 211, 213, 211, 213, 210, 207, 209, 211, 209, 209, 206, 211, 206, 207, 208, 205, 211, 209, 205, 211, 214, 212, 211, 211, 211, 212, 211, 212, 211, 211, 209, 214, 212, 212, 208, 204, 206, 207, 207, 205, 205, 208, 207, 207, 210, 208, 206, 210, 206, 201, 197, 202, 192, 138, 192, 190, 187, 191, 116, 189, 195, 193, 192, 191, 194, 194, 192, 198, 198, 196, 197, 199, 202, 201, 198, 197, 197, 200, 200, 197, 199, 197, 199, 199, 200, 202, 206, 202, 202, 204, 202, 202, 200, 198, 203, 202, 205, 203, 205, 205, 209, 207, 206, 205, 207, 206, 208, 207, 207, 208, 206, 204, 206, 204, 208, 206, 207, 209, 207, 210, 211, 214, 215, 212, 210, 208, 213, 213, 211, 209, 211, 208, 209, 213, 211, 212, 212, 212, 214, 209, 211, 212, 214, 216, 213, 211, 214, 211, 214, 216, 215, 213, 215, 213, 213, 213, 215, 215, 217, 213, 215, 213, 212, 214, 214, 218, 216, 216, 214, 214, 215, 211, 213, 209, 210, 214, 216, 214, 216, 214, 212, 211, 212, 212, 212, 215, 211, 213, 216, 215, 218, 216, 216, 216, 215, 214, 213, 216, 213, 213, 216, 216, 216, 217, 215, 214, 215, 214, 213, 216, 217, 215, 214, 210, 212, 212, 214, 213, 210, 212, 212, 213, 218, 214, 210, 216, 213, 213, 212, 209, 215, 213, 213, 215, 210, 209, 214, 209, 210, 204, 205, 206, 212, 210, 210, 211, 209, 205, 212, 212, 210, 207, 210, 211, 215, 212, 213, 212, 214, 214, 209, 207, 211, 210, 209, 212, 208, 209, 213, 207, 210, 211, 210, 209, 212, 214, 215, 215, 211, 210, 212, 212, 213, 214, 213, 211, 211, 209, 210, 209, 207, 210, 209, 213, 207, 207, 208, 207, 209, 207, 208, 211, 208, 209, 211, 205, 202, 198, 191, 145, 195, 195, 189, 196, 116, 192, 193, 196, 193, 197, 198, 197, 198, 197, 199, 194, 197, 199, 205, 199, 200, 201, 202, 201, 201, 198, 201, 201, 199, 199, 200, 202, 201, 203, 202, 208, 203, 205, 203, 202, 204, 201, 206, 203, 208, 206, 206, 208, 209, 208, 210, 210, 209, 203, 209, 207, 207, 207, 206, 207, 209, 204, 210, 208, 212, 211, 212, 213, 213, 213, 210, 209, 210, 210, 212, 211, 207, 210, 211, 214, 213, 209, 209, 212, 217, 211, 212, 213, 215, 216, 212, 208, 212, 210, 212, 214, 216, 212, 211, 214, 213, 212, 213, 212, 212, 211, 214, 214, 210, 214, 218, 217, 216, 217, 217, 214, 212, 210, 212, 209, 212, 213, 215, 213, 215, 213, 213, 211, 210, 211, 213, 212, 212, 214, 217, 214, 217, 216, 216, 215, 213, 213, 215, 215, 218, 214, 216, 214, 214, 215, 219, 218, 215, 216, 217, 215, 219, 214, 214, 213, 215, 212, 213, 214, 214, 216, 215, 215, 220, 217, 215, 214, 217, 214, 211, 211, 213, 212, 215, 213, 210, 208, 212, 210, 211, 205, 204, 208, 212, 212, 208, 212, 212, 209, 212, 211, 208, 208, 210, 210, 213, 213, 215, 214, 216, 213, 210, 210, 209, 211, 208, 211, 209, 207, 211, 209, 210, 207, 208, 210, 214, 214, 218, 215, 213, 215, 215, 215, 215, 215, 213, 210, 211, 213, 215, 210, 205, 210, 209, 213, 208, 208, 211, 211, 213, 215, 209, 208, 209, 207, 210, 207, 203, 200, 198, 150, 194, 195, 189, 195, 130, 192, 199, 192, 192, 197, 195, 195, 197, 194, 198, 196, 197, 201, 197, 201, 201, 196, 201, 203, 202, 201, 198, 197, 196, 198, 203, 205, 206, 207, 204, 204, 205, 205, 204, 205, 206, 204, 206, 203, 207, 209, 208, 206, 208, 208, 209, 209, 209, 205, 208, 211, 205, 210, 209, 209, 210, 208, 211, 210, 211, 209, 212, 212, 214, 213, 208, 212, 209, 212, 212, 216, 210, 215, 214, 213, 212, 210, 212, 213, 211, 210, 210, 212, 213, 211, 204, 210, 212, 213, 214, 213, 213, 213, 211, 216, 213, 214, 214, 213, 213, 212, 214, 211, 212, 216, 215, 219, 217, 218, 218, 214, 214, 211, 212, 213, 213, 212, 215, 213, 214, 211, 212, 214, 212, 213, 212, 211, 214, 216, 218, 216, 217, 216, 214, 215, 215, 217, 217, 217, 215, 216, 216, 217, 216, 217, 219, 217, 215, 214, 215, 215, 217, 216, 215, 218, 215, 214, 213, 217, 218, 216, 216, 217, 215, 217, 214, 216, 217, 217, 214, 212, 213, 214, 216, 215, 212, 213, 211, 213, 212, 207, 206, 212, 213, 212, 212, 213, 211, 211, 213, 214, 211, 209, 209, 213, 216, 216, 213, 213, 216, 213, 212, 211, 208, 214, 208, 211, 211, 209, 214, 208, 214, 215, 210, 213, 217, 214, 214, 215, 213, 214, 216, 214, 216, 214, 213, 217, 214, 214, 210, 211, 209, 210, 210, 214, 211, 210, 211, 209, 212, 217, 209, 212, 209, 207, 207, 207, 206, 202, 198, 161, 195, 195, 189, 192, 115, 195, 194, 194, 196, 201, 196, 200, 195, 195, 199, 200, 198, 202, 201, 199, 200, 200, 202, 200, 201, 204, 201, 200, 200, 200, 203, 207, 206, 206, 205, 201, 207, 207, 206, 206, 207, 202, 202, 203, 204, 206, 208, 209, 209, 209, 210, 213, 209, 205, 208, 207, 204, 208, 209, 208, 212, 211, 212, 213, 210, 211, 212, 213, 214, 214, 210, 211, 212, 214, 214, 216, 212, 214, 212, 211, 211, 210, 212, 212, 213, 213, 210, 209, 213, 216, 209, 213, 216, 215, 213, 216, 214, 209, 209, 214, 216, 212, 213, 212, 214, 215, 214, 212, 215, 215, 214, 218, 217, 216, 217, 217, 214, 209, 213, 214, 212, 210, 213, 212, 212, 211, 213, 215, 211, 213, 216, 214, 215, 216, 219, 217, 216, 212, 217, 214, 216, 216, 216, 217, 217, 218, 215, 214, 217, 218, 217, 218, 217, 218, 215, 218, 217, 216, 215, 215, 214, 216, 218, 219, 219, 218, 215, 217, 215, 214, 213, 215, 218, 215, 216, 215, 214, 216, 218, 218, 211, 213, 216, 218, 216, 213, 213, 209, 215, 213, 215, 212, 215, 213, 216, 214, 212, 211, 213, 212, 213, 215, 213, 216, 215, 211, 214, 210, 209, 211, 213, 213, 212, 213, 216, 214, 212, 213, 215, 214, 216, 216, 219, 214, 212, 215, 213, 215, 215, 211, 214, 215, 215, 214, 211, 213, 208, 208, 212, 207, 214, 209, 208, 211, 208, 207, 209, 210, 206, 208, 207, 206, 211, 204, 198, 175, 198, 190, 189, 191, 124, 192, 197, 195, 194, 199, 200, 197, 194, 195, 197, 201, 197, 199, 200, 198, 202, 198, 205, 203, 205, 203, 203, 204, 203, 201, 202, 203, 202, 203, 205, 205, 204, 207, 204, 206, 205, 204, 204, 204, 206, 205, 211, 207, 207, 210, 212, 213, 209, 210, 209, 211, 208, 208, 208, 206, 209, 209, 210, 209, 209, 210, 212, 211, 210, 212, 210, 210, 209, 214, 213, 212, 213, 211, 214, 213, 213, 209, 209, 213, 214, 213, 215, 212, 215, 216, 215, 216, 214, 214, 215, 213, 215, 213, 214, 215, 214, 217, 216, 217, 217, 214, 216, 212, 212, 214, 213, 215, 214, 216, 214, 214, 218, 211, 214, 214, 214, 212, 213, 212, 210, 213, 215, 211, 214, 215, 214, 216, 215, 216, 219, 216, 216, 215, 215, 216, 217, 220, 216, 215, 220, 220, 216, 216, 218, 217, 218, 219, 217, 217, 217, 218, 220, 217, 219, 216, 215, 218, 218, 219, 219, 218, 220, 218, 214, 213, 213, 215, 218, 220, 217, 214, 212, 210, 216, 216, 210, 214, 214, 216, 214, 214, 214, 212, 212, 213, 215, 212, 213, 216, 214, 212, 209, 209, 213, 215, 212, 216, 209, 216, 216, 213, 213, 213, 211, 212, 210, 212, 213, 210, 214, 214, 213, 216, 217, 214, 215, 214, 217, 213, 212, 211, 212, 215, 213, 213, 213, 213, 212, 211, 210, 212, 211, 208, 212, 213, 213, 212, 212, 210, 207, 209, 210, 207, 207, 210, 209, 209, 206, 205, 196, 166, 195, 190, 191, 196, 132, 195, 197, 198, 197, 197, 198, 198, 197, 196, 197, 198, 203, 202, 201, 199, 199, 200, 200, 203, 200, 199, 200, 200, 200, 200, 206, 203, 202, 202, 206, 209, 207, 205, 206, 205, 205, 205, 207, 209, 209, 209, 210, 208, 209, 213, 214, 209, 212, 208, 210, 211, 212, 211, 212, 209, 208, 212, 213, 213, 212, 211, 209, 208, 210, 209, 208, 211, 212, 214, 212, 215, 215, 212, 214, 213, 212, 210, 210, 214, 212, 213, 212, 215, 214, 216, 214, 214, 214, 217, 219, 216, 215, 213, 213, 213, 216, 216, 213, 217, 216, 217, 218, 214, 214, 216, 214, 216, 218, 218, 216, 214, 213, 215, 212, 213, 211, 210, 212, 210, 210, 214, 213, 214, 216, 214, 213, 216, 218, 218, 216, 216, 216, 215, 217, 217, 218, 218, 220, 219, 221, 222, 220, 218, 217, 218, 219, 218, 217, 216, 217, 216, 220, 218, 215, 215, 218, 217, 218, 218, 219, 217, 217, 216, 216, 214, 215, 212, 217, 215, 215, 212, 211, 212, 215, 214, 215, 216, 219, 214, 217, 214, 212, 215, 216, 212, 210, 216, 214, 216, 214, 212, 212, 213, 211, 219, 212, 213, 212, 217, 216, 216, 213, 216, 213, 211, 213, 217, 216, 211, 213, 214, 213, 214, 217, 218, 216, 214, 215, 217, 212, 211, 214, 212, 215, 214, 216, 214, 214, 210, 209, 212, 212, 214, 214, 214, 213, 213, 214, 210, 211, 208, 210, 207, 210, 209, 212, 211, 206, 207, 199, 156, 193, 191, 193, 198, 134, 190, 196, 198, 193, 198, 198, 199, 199, 200, 200, 200, 200, 201, 203, 202, 199, 201, 202, 204, 199, 202, 202, 202, 199, 204, 206, 205, 203, 206, 204, 207, 204, 206, 205, 205, 205, 205, 207, 207, 214, 210, 212, 208, 210, 213, 211, 210, 214, 210, 212, 212, 212, 211, 207, 208, 210, 208, 215, 213, 211, 213, 213, 213, 211, 211, 211, 209, 214, 215, 214, 214, 216, 214, 214, 213, 212, 211, 212, 215, 214, 212, 208, 215, 215, 216, 219, 214, 216, 216, 218, 219, 216, 215, 214, 218, 217, 218, 218, 220, 218, 218, 216, 217, 216, 213, 216, 218, 218, 216, 217, 214, 217, 217, 215, 214, 212, 210, 215, 214, 216, 215, 215, 215, 216, 214, 210, 216, 217, 216, 216, 216, 216, 214, 215, 216, 221, 219, 219, 218, 223, 221, 223, 219, 217, 219, 218, 219, 216, 217, 216, 221, 220, 217, 213, 216, 220, 218, 217, 216, 217, 218, 220, 220, 218, 215, 216, 216, 218, 218, 218, 213, 212, 213, 216, 216, 216, 210, 214, 217, 218, 213, 210, 214, 213, 213, 215, 215, 215, 216, 215, 216, 216, 217, 213, 216, 211, 213, 213, 212, 215, 214, 215, 215, 217, 216, 212, 212, 217, 214, 214, 214, 212, 215, 219, 216, 215, 218, 219, 216, 215, 214, 213, 213, 214, 218, 215, 215, 212, 212, 215, 215, 217, 214, 217, 214, 212, 214, 212, 211, 213, 208, 209, 208, 209, 209, 211, 210, 208, 205, 197, 145, 195, 195, 192, 197, 121, 194, 194, 193, 198, 196, 198, 201, 200, 196, 197, 193, 195, 203, 199, 203, 199, 201, 203, 204, 203, 204, 201, 201, 201, 203, 206, 201, 203, 205, 205, 209, 204, 208, 205, 206, 205, 207, 206, 210, 210, 211, 213, 211, 210, 213, 213, 213, 213, 208, 212, 212, 211, 212, 211, 206, 212, 213, 218, 208, 211, 212, 216, 215, 210, 213, 214, 214, 212, 215, 214, 213, 212, 214, 212, 212, 209, 213, 208, 214, 211, 213, 214, 214, 215, 219, 217, 214, 218, 217, 218, 217, 217, 216, 213, 215, 216, 215, 217, 217, 215, 216, 217, 217, 219, 216, 219, 218, 218, 216, 213, 218, 215, 215, 215, 213, 212, 216, 215, 216, 213, 216, 216, 218, 215, 215, 215, 217, 218, 217, 217, 215, 216, 213, 216, 218, 220, 219, 218, 218, 221, 221, 221, 219, 221, 220, 218, 220, 216, 218, 218, 218, 218, 218, 217, 216, 219, 218, 219, 219, 219, 216, 218, 217, 215, 216, 221, 216, 219, 218, 218, 214, 210, 216, 214, 217, 213, 212, 215, 217, 214, 213, 213, 215, 216, 214, 215, 214, 212, 219, 215, 213, 215, 218, 218, 216, 210, 217, 215, 214, 213, 213, 214, 215, 215, 216, 218, 214, 214, 214, 212, 214, 219, 216, 219, 218, 216, 217, 217, 216, 215, 214, 213, 213, 217, 216, 211, 214, 216, 217, 216, 215, 216, 212, 217, 213, 215, 215, 211, 213, 213, 212, 209, 211, 209, 210, 212, 211, 208, 205, 197, 145, 196, 194, 192, 198, 117, 195, 199, 197, 198, 198, 198, 201, 197, 196, 195, 197, 198, 202, 201, 202, 200, 198, 206, 203, 205, 206, 203, 204, 204, 203, 206, 204, 204, 204, 206, 206, 207, 207, 205, 207, 206, 206, 211, 210, 212, 211, 213, 211, 210, 211, 210, 211, 212, 208, 209, 216, 210, 207, 211, 210, 210, 213, 216, 213, 213, 213, 216, 218, 215, 213, 212, 214, 215, 214, 215, 212, 210, 213, 216, 212, 212, 212, 210, 212, 213, 213, 215, 215, 217, 217, 217, 215, 217, 213, 215, 220, 218, 216, 215, 214, 216, 219, 214, 217, 219, 218, 217, 217, 217, 217, 216, 216, 217, 216, 218, 218, 217, 217, 215, 216, 215, 216, 215, 216, 214, 219, 217, 216, 217, 220, 217, 218, 217, 216, 215, 215, 217, 213, 218, 221, 220, 218, 220, 220, 220, 221, 220, 218, 219, 218, 218, 217, 217, 217, 221, 221, 218, 218, 216, 218, 219, 219, 220, 216, 216, 217, 216, 217, 216, 218, 219, 219, 219, 220, 217, 216, 216, 217, 218, 214, 210, 212, 213, 216, 214, 214, 217, 214, 217, 216, 216, 216, 217, 215, 219, 215, 215, 214, 215, 217, 215, 213, 216, 214, 214, 215, 212, 216, 215, 215, 218, 217, 217, 213, 213, 212, 213, 214, 218, 217, 215, 219, 218, 217, 215, 217, 216, 216, 214, 216, 213, 214, 217, 216, 216, 215, 215, 215, 214, 217, 218, 215, 213, 213, 213, 214, 209, 210, 210, 213, 214, 211, 209, 205, 199, 150, 199, 197, 194, 199, 126, 195, 201, 200, 195, 200, 196, 201, 203, 196, 201, 198, 195, 201, 198, 199, 204, 203, 208, 204, 205, 206, 204, 205, 205, 202, 205, 205, 208, 204, 209, 207, 207, 207, 206, 206, 208, 206, 206, 208, 210, 210, 211, 211, 209, 208, 211, 210, 211, 209, 212, 213, 209, 213, 211, 213, 212, 213, 215, 212, 212, 211, 215, 214, 211, 211, 212, 215, 217, 213, 215, 214, 209, 214, 214, 215, 213, 212, 211, 215, 211, 216, 214, 216, 216, 218, 216, 217, 215, 214, 218, 220, 216, 213, 217, 218, 213, 218, 218, 216, 220, 219, 220, 219, 217, 214, 217, 218, 217, 216, 217, 216, 218, 219, 217, 217, 216, 217, 215, 218, 218, 217, 214, 213, 215, 217, 217, 215, 215, 216, 219, 216, 221, 216, 217, 220, 223, 219, 220, 220, 221, 222, 221, 220, 220, 218, 219, 221, 219, 216, 220, 218, 219, 220, 217, 220, 219, 219, 218, 215, 216, 216, 216, 216, 214, 219, 219, 218, 221, 220, 217, 216, 214, 217, 216, 211, 213, 214, 217, 218, 213, 215, 213, 214, 218, 217, 217, 216, 218, 217, 217, 216, 218, 213, 216, 217, 216, 217, 215, 217, 217, 216, 216, 217, 217, 217, 217, 219, 216, 214, 212, 211, 213, 215, 215, 216, 214, 218, 217, 216, 217, 214, 216, 217, 217, 215, 218, 215, 217, 216, 218, 215, 213, 215, 214, 217, 217, 217, 213, 214, 212, 214, 211, 212, 211, 212, 216, 214, 207, 205, 201, 159, 198, 193, 192, 201, 124, 192, 199, 197, 196, 196, 200, 200, 200, 196, 198, 195, 197, 207, 204, 207, 201, 206, 207, 205, 210, 207, 210, 207, 210, 206, 204, 208, 206, 205, 207, 207, 208, 206, 208, 205, 206, 206, 207, 211, 210, 212, 213, 211, 210, 212, 214, 214, 213, 211, 214, 213, 210, 213, 211, 214, 215, 214, 214, 214, 215, 212, 214, 213, 213, 214, 217, 214, 216, 214, 212, 212, 213, 214, 218, 219, 212, 212, 211, 215, 214, 213, 216, 212, 216, 220, 220, 219, 216, 216, 218, 221, 216, 213, 215, 216, 216, 220, 221, 219, 218, 220, 218, 217, 218, 214, 217, 218, 216, 221, 216, 215, 217, 216, 215, 217, 216, 217, 216, 216, 215, 216, 218, 215, 215, 218, 216, 217, 216, 215, 217, 217, 217, 217, 218, 222, 221, 218, 222, 221, 221, 221, 222, 222, 220, 220, 220, 219, 221, 217, 218, 221, 220, 217, 217, 218, 217, 220, 218, 217, 218, 215, 221, 221, 219, 220, 217, 221, 221, 218, 214, 216, 220, 216, 218, 215, 215, 213, 218, 217, 215, 215, 214, 212, 216, 216, 217, 219, 219, 219, 221, 218, 216, 215, 215, 218, 218, 218, 216, 215, 216, 217, 218, 215, 216, 217, 219, 219, 214, 214, 215, 216, 218, 217, 218, 217, 219, 221, 219, 215, 216, 215, 218, 217, 217, 216, 215, 213, 214, 217, 216, 214, 213, 213, 215, 214, 212, 216, 213, 210, 212, 216, 208, 210, 211, 215, 216, 213, 211, 208, 198, 155, 202, 193, 195, 196, 117, 193, 201, 198, 196, 196, 202, 198, 201, 199, 197, 198, 197, 199, 206, 205, 209, 206, 209, 208, 209, 209, 209, 206, 210, 202, 203, 208, 203, 204, 206, 206, 205, 205, 206, 208, 209, 206, 211, 212, 215, 214, 213, 211, 210, 213, 216, 213, 211, 211, 214, 215, 213, 213, 216, 217, 217, 215, 218, 214, 216, 212, 213, 216, 214, 216, 216, 216, 214, 216, 210, 212, 212, 213, 217, 217, 215, 213, 215, 216, 213, 211, 214, 215, 216, 217, 218, 217, 214, 215, 221, 217, 217, 217, 214, 218, 217, 218, 220, 216, 219, 220, 219, 217, 216, 217, 219, 218, 218, 220, 219, 216, 220, 219, 218, 220, 219, 216, 217, 216, 215, 216, 219, 218, 218, 219, 216, 217, 212, 218, 219, 215, 216, 217, 223, 223, 223, 221, 222, 222, 224, 221, 221, 223, 222, 222, 218, 219, 217, 216, 218, 222, 218, 218, 217, 221, 219, 220, 218, 217, 214, 221, 221, 221, 222, 219, 221, 223, 222, 218, 218, 217, 218, 219, 218, 215, 214, 215, 215, 218, 218, 215, 216, 216, 218, 219, 218, 218, 218, 219, 219, 219, 217, 219, 215, 216, 219, 217, 222, 215, 217, 219, 219, 218, 216, 216, 221, 219, 218, 214, 216, 216, 218, 217, 217, 216, 221, 220, 220, 216, 216, 213, 216, 220, 216, 217, 219, 218, 215, 218, 219, 217, 217, 214, 217, 217, 215, 215, 214, 213, 213, 213, 213, 209, 212, 215, 213, 215, 211, 204, 198, 159, 202, 196, 192, 199, 103, 189, 198, 197, 197, 198, 195, 201, 199, 198, 195, 198, 197, 199, 205, 202, 205, 207, 208, 207, 208, 206, 205, 204, 207, 202, 202, 203, 205, 207, 205, 208, 208, 205, 204, 210, 212, 209, 213, 210, 212, 213, 210, 211, 207, 214, 214, 213, 214, 213, 217, 216, 217, 215, 214, 215, 218, 217, 219, 216, 212, 213, 214, 217, 216, 214, 218, 219, 216, 214, 214, 210, 212, 214, 215, 214, 215, 215, 215, 215, 215, 214, 217, 214, 217, 216, 219, 221, 217, 217, 220, 220, 216, 214, 217, 220, 220, 218, 219, 216, 220, 219, 218, 218, 216, 218, 220, 217, 219, 217, 217, 218, 218, 218, 219, 218, 218, 215, 215, 216, 217, 216, 217, 219, 215, 218, 215, 214, 216, 219, 219, 218, 219, 219, 222, 222, 222, 223, 222, 221, 223, 220, 219, 220, 221, 220, 218, 218, 218, 218, 219, 223, 223, 218, 218, 221, 220, 221, 218, 216, 218, 219, 220, 219, 218, 218, 219, 224, 223, 220, 217, 216, 217, 217, 217, 217, 214, 215, 216, 216, 215, 217, 216, 219, 217, 218, 216, 216, 220, 218, 219, 216, 212, 216, 216, 219, 217, 218, 215, 214, 218, 216, 216, 219, 216, 215, 218, 216, 215, 220, 216, 216, 218, 216, 217, 217, 217, 219, 219, 218, 218, 215, 216, 219, 221, 217, 216, 214, 218, 216, 216, 215, 215, 216, 212, 214, 214, 212, 215, 215, 214, 216, 211, 213, 209, 213, 216, 216, 212, 207, 196, 151, 199, 196, 195, 198, 115, 193, 199, 194, 194, 196, 198, 202, 199, 197, 198, 201, 201, 203, 203, 205, 206, 205, 206, 205, 208, 203, 207, 208, 206, 205, 210, 205, 205, 204, 207, 210, 209, 209, 205, 211, 209, 210, 210, 214, 212, 212, 209, 208, 208, 214, 215, 212, 214, 214, 214, 212, 216, 214, 218, 216, 216, 216, 219, 212, 212, 215, 216, 217, 214, 217, 219, 221, 219, 216, 218, 212, 209, 213, 214, 215, 216, 214, 214, 215, 216, 217, 216, 215, 218, 218, 218, 220, 221, 216, 221, 218, 218, 217, 214, 219, 219, 220, 219, 218, 218, 220, 218, 220, 217, 215, 217, 219, 218, 218, 218, 218, 218, 218, 221, 219, 218, 215, 218, 215, 215, 218, 218, 217, 220, 217, 218, 217, 218, 218, 216, 220, 219, 218, 220, 221, 225, 221, 222, 221, 222, 221, 220, 220, 222, 220, 222, 221, 217, 219, 222, 220, 221, 223, 223, 218, 220, 223, 221, 216, 218, 218, 220, 222, 219, 220, 221, 224, 223, 223, 221, 217, 218, 218, 218, 217, 211, 216, 216, 216, 215, 213, 218, 219, 220, 220, 216, 216, 218, 219, 219, 218, 217, 217, 216, 218, 217, 222, 218, 217, 220, 218, 218, 218, 217, 216, 218, 216, 214, 219, 215, 215, 218, 219, 216, 217, 217, 219, 219, 217, 218, 217, 217, 220, 221, 220, 217, 217, 220, 215, 217, 217, 213, 213, 213, 218, 217, 215, 212, 214, 215, 217, 211, 214, 208, 215, 213, 213, 213, 209, 203, 156, 198, 198, 195, 198, 103, 192, 194, 196, 192, 201, 199, 202, 198, 198, 203, 197, 202, 202, 202, 206, 208, 207, 209, 207, 204, 205, 206, 206, 211, 209, 213, 208, 206, 207, 209, 209, 207, 208, 209, 211, 213, 211, 211, 209, 211, 212, 209, 210, 209, 213, 216, 211, 214, 213, 218, 214, 217, 215, 217, 214, 217, 216, 217, 212, 216, 215, 218, 216, 215, 217, 217, 219, 217, 220, 215, 217, 213, 217, 215, 216, 216, 217, 216, 217, 217, 216, 216, 215, 219, 219, 219, 220, 219, 216, 219, 220, 218, 217, 217, 219, 220, 219, 220, 219, 219, 222, 219, 219, 215, 216, 218, 216, 220, 219, 221, 218, 219, 219, 219, 216, 217, 216, 218, 218, 218, 215, 219, 216, 218, 216, 218, 219, 219, 220, 219, 220, 221, 221, 218, 221, 223, 219, 221, 223, 223, 220, 221, 222, 222, 223, 222, 218, 218, 218, 222, 222, 223, 223, 222, 220, 220, 222, 221, 218, 218, 218, 220, 223, 222, 219, 222, 223, 221, 224, 220, 218, 221, 219, 219, 219, 214, 216, 216, 217, 216, 213, 221, 216, 217, 215, 217, 218, 218, 218, 218, 219, 218, 216, 220, 218, 221, 219, 220, 219, 220, 218, 218, 221, 216, 216, 216, 215, 219, 219, 218, 215, 216, 217, 219, 215, 218, 217, 218, 219, 217, 216, 216, 221, 217, 222, 218, 218, 220, 216, 218, 213, 214, 210, 219, 216, 213, 217, 215, 217, 216, 215, 214, 213, 213, 215, 217, 216, 210, 210, 202, 154, 202, 194, 197, 197, 91, 192, 197, 196, 198, 200, 198, 200, 202, 201, 198, 201, 202, 204, 205, 206, 208, 209, 208, 208, 206, 205, 208, 207, 211, 209, 211, 208, 211, 209, 210, 208, 206, 209, 212, 210, 212, 212, 214, 210, 212, 213, 211, 209, 212, 212, 216, 216, 217, 216, 216, 215, 217, 217, 213, 217, 219, 216, 218, 216, 216, 217, 216, 219, 214, 216, 216, 217, 217, 216, 216, 218, 215, 216, 218, 217, 217, 219, 216, 220, 216, 217, 218, 217, 219, 216, 219, 220, 218, 216, 218, 219, 221, 218, 218, 219, 220, 217, 222, 222, 220, 222, 220, 218, 215, 216, 221, 220, 223, 223, 220, 217, 220, 221, 221, 218, 216, 215, 221, 219, 219, 214, 220, 216, 216, 218, 218, 218, 217, 218, 220, 219, 222, 220, 222, 220, 223, 220, 222, 224, 223, 222, 224, 221, 221, 223, 221, 221, 219, 221, 220, 223, 222, 223, 219, 222, 224, 225, 222, 219, 222, 220, 218, 223, 221, 219, 218, 221, 221, 220, 219, 219, 221, 220, 219, 220, 216, 217, 220, 218, 218, 217, 221, 218, 220, 213, 219, 218, 219, 218, 217, 219, 213, 217, 220, 218, 220, 220, 221, 221, 219, 216, 221, 221, 217, 214, 216, 215, 218, 219, 220, 215, 218, 219, 221, 216, 216, 217, 217, 220, 217, 216, 219, 220, 223, 221, 219, 218, 217, 215, 214, 213, 211, 213, 215, 218, 217, 219, 217, 218, 217, 217, 212, 213, 214, 212, 216, 214, 213, 208, 201, 156, 200, 198, 195, 198, 89, 190, 198, 196, 196, 198, 201, 200, 201, 203, 200, 203, 207, 208, 206, 207, 205, 206, 211, 203, 210, 210, 210, 210, 211, 210, 209, 209, 210, 211, 210, 210, 207, 210, 212, 211, 212, 214, 212, 212, 211, 211, 213, 213, 212, 213, 213, 217, 217, 217, 216, 216, 218, 216, 214, 218, 217, 217, 219, 217, 216, 217, 218, 219, 215, 218, 215, 216, 216, 220, 216, 217, 216, 216, 220, 217, 219, 218, 218, 219, 216, 218, 216, 217, 218, 217, 219, 217, 218, 216, 218, 220, 217, 220, 218, 219, 220, 221, 221, 222, 219, 219, 219, 220, 216, 220, 220, 221, 218, 221, 221, 221, 221, 223, 220, 218, 217, 217, 221, 220, 219, 217, 218, 217, 218, 219, 217, 219, 218, 218, 218, 218, 221, 222, 220, 222, 222, 224, 222, 224, 223, 222, 224, 220, 219, 223, 219, 220, 221, 219, 220, 224, 223, 221, 219, 223, 224, 222, 222, 220, 219, 220, 218, 222, 221, 219, 219, 220, 221, 222, 215, 220, 220, 222, 220, 219, 217, 221, 220, 219, 219, 217, 219, 216, 220, 218, 222, 218, 221, 220, 218, 216, 218, 217, 219, 220, 219, 219, 220, 220, 219, 220, 216, 217, 216, 216, 219, 218, 217, 219, 220, 216, 218, 221, 219, 217, 216, 220, 221, 222, 220, 218, 220, 224, 222, 221, 220, 217, 217, 218, 218, 214, 211, 216, 218, 217, 214, 219, 216, 220, 216, 218, 215, 215, 215, 213, 218, 217, 214, 209, 202, 152, 203, 201, 198, 200, 91, 193, 198, 195, 197, 196, 195, 201, 197, 202, 201, 203, 202, 206, 206, 209, 212, 210, 211, 207, 209, 209, 205, 210, 207, 211, 210, 212, 209, 210, 210, 209, 209, 212, 213, 214, 212, 215, 210, 212, 212, 212, 215, 213, 214, 215, 213, 216, 218, 214, 217, 218, 218, 217, 215, 217, 218, 218, 219, 217, 217, 218, 217, 223, 216, 218, 218, 218, 220, 220, 218, 217, 215, 216, 219, 213, 216, 216, 220, 219, 217, 220, 218, 218, 218, 218, 219, 217, 218, 217, 220, 222, 221, 219, 219, 220, 220, 223, 219, 221, 219, 221, 223, 220, 218, 219, 222, 221, 220, 222, 220, 223, 222, 222, 219, 218, 219, 219, 222, 219, 220, 219, 218, 219, 219, 219, 218, 219, 219, 219, 217, 219, 222, 222, 223, 224, 223, 223, 224, 223, 225, 222, 222, 220, 219, 221, 223, 220, 220, 219, 221, 223, 223, 223, 222, 222, 222, 224, 222, 221, 221, 221, 220, 224, 221, 220, 218, 221, 222, 221, 217, 218, 220, 224, 219, 218, 217, 219, 223, 220, 219, 220, 217, 216, 220, 221, 219, 220, 221, 219, 219, 217, 218, 220, 215, 220, 218, 217, 221, 222, 221, 218, 218, 215, 215, 217, 218, 218, 218, 217, 219, 217, 220, 221, 218, 220, 221, 219, 222, 224, 218, 217, 218, 220, 221, 221, 221, 220, 222, 218, 220, 215, 213, 218, 220, 219, 219, 218, 215, 218, 216, 220, 218, 215, 215, 214, 220, 216, 215, 214, 206, 155, 200, 199, 195, 199, 109, 197, 202, 197, 197, 195, 199, 203, 202, 204, 200, 203, 208, 207, 207, 206, 210, 211, 210, 207, 207, 205, 206, 208, 215, 211, 210, 210, 212, 211, 208, 208, 208, 212, 209, 215, 212, 213, 212, 210, 215, 211, 212, 212, 213, 212, 217, 216, 216, 217, 215, 219, 217, 216, 215, 216, 216, 217, 219, 218, 219, 218, 219, 221, 217, 217, 219, 218, 221, 220, 218, 218, 218, 218, 218, 216, 216, 217, 220, 221, 220, 221, 219, 215, 217, 220, 216, 219, 217, 217, 221, 220, 221, 219, 221, 220, 221, 222, 219, 221, 221, 223, 224, 223, 223, 221, 221, 222, 221, 222, 222, 220, 223, 221, 220, 218, 219, 219, 223, 220, 219, 220, 218, 221, 219, 221, 218, 220, 223, 222, 221, 218, 221, 222, 220, 222, 225, 221, 224, 223, 222, 224, 222, 221, 221, 221, 219, 220, 222, 221, 220, 222, 223, 221, 224, 221, 223, 223, 224, 220, 222, 221, 221, 225, 222, 220, 217, 220, 221, 223, 219, 219, 222, 223, 222, 218, 221, 219, 219, 218, 219, 221, 219, 220, 219, 221, 221, 220, 219, 219, 219, 221, 218, 219, 217, 221, 222, 220, 222, 220, 219, 218, 220, 214, 218, 216, 220, 221, 220, 217, 219, 217, 221, 220, 218, 221, 219, 222, 224, 221, 218, 216, 219, 219, 222, 219, 219, 221, 222, 221, 221, 217, 217, 219, 219, 217, 218, 218, 217, 219, 217, 222, 216, 217, 217, 219, 218, 215, 220, 215, 206, 175, 203, 197, 199, 200, 97, 198, 201, 198, 198, 195, 200, 200, 203, 202, 203, 206, 209, 205, 207, 206, 204, 209, 206, 211, 208, 206, 208, 208, 213, 215, 209, 212, 208, 214, 212, 211, 212, 207, 211, 212, 212, 211, 212, 212, 213, 213, 214, 218, 216, 216, 213, 217, 214, 217, 219, 218, 217, 218, 217, 216, 213, 216, 218, 218, 219, 218, 220, 220, 219, 219, 220, 218, 221, 221, 220, 220, 220, 220, 220, 216, 217, 219, 218, 221, 220, 220, 219, 217, 217, 219, 218, 222, 222, 223, 224, 222, 223, 221, 217, 220, 222, 222, 223, 220, 221, 223, 225, 223, 223, 223, 221, 222, 221, 220, 222, 220, 224, 224, 223, 221, 218, 218, 222, 222, 220, 219, 220, 217, 222, 223, 217, 217, 219, 221, 221, 220, 216, 222, 222, 224, 225, 222, 224, 223, 224, 224, 222, 217, 222, 223, 221, 222, 220, 222, 222, 224, 225, 220, 224, 221, 224, 224, 224, 221, 219, 221, 224, 222, 222, 218, 218, 223, 223, 224, 221, 220, 222, 222, 222, 219, 217, 217, 220, 219, 223, 218, 220, 221, 221, 222, 222, 218, 222, 221, 220, 222, 219, 218, 219, 224, 223, 220, 222, 222, 221, 221, 219, 215, 215, 218, 224, 220, 220, 218, 218, 219, 223, 223, 220, 221, 219, 225, 222, 223, 217, 222, 221, 221, 220, 220, 221, 219, 220, 221, 222, 221, 219, 219, 220, 217, 217, 218, 217, 217, 218, 217, 214, 218, 219, 219, 218, 218, 221, 215, 206, 189, 206, 199, 196, 202, 98, 195, 198, 200, 195, 197, 198, 200, 201, 200, 203, 202, 206, 206, 207, 206, 207, 208, 208, 206, 209, 207, 207, 208, 211, 212, 208, 211, 207, 213, 212, 209, 209, 211, 213, 214, 210, 213, 211, 213, 216, 215, 218, 219, 214, 216, 217, 218, 216, 215, 219, 215, 218, 220, 220, 216, 222, 218, 219, 219, 217, 219, 221, 222, 218, 217, 221, 218, 223, 220, 222, 218, 219, 217, 220, 220, 220, 218, 220, 220, 220, 218, 220, 217, 222, 220, 221, 221, 220, 222, 224, 223, 222, 220, 220, 220, 223, 224, 221, 221, 222, 225, 222, 222, 222, 223, 223, 224, 221, 220, 224, 221, 225, 224, 224, 219, 221, 220, 223, 222, 220, 219, 219, 220, 221, 221, 220, 219, 219, 222, 220, 218, 221, 223, 222, 225, 226, 225, 223, 223, 222, 225, 223, 222, 225, 223, 221, 224, 219, 223, 221, 226, 225, 223, 222, 222, 223, 226, 224, 223, 222, 222, 225, 221, 222, 223, 220, 222, 221, 220, 219, 220, 221, 221, 222, 221, 217, 217, 223, 221, 223, 220, 221, 222, 222, 219, 219, 218, 218, 221, 221, 221, 222, 219, 220, 224, 222, 220, 220, 221, 220, 218, 219, 218, 220, 220, 224, 222, 222, 219, 220, 220, 223, 221, 222, 221, 219, 222, 220, 224, 222, 221, 222, 219, 223, 222, 221, 220, 220, 224, 223, 223, 224, 220, 222, 221, 217, 221, 217, 220, 219, 215, 214, 218, 217, 219, 222, 220, 221, 214, 212, 189, 201, 200, 201, 203, 99, 198, 204, 205, 197, 199, 200, 202, 203, 202, 207, 208, 207, 207, 205, 199, 205, 208, 205, 205, 209, 207, 209, 211, 211, 210, 208, 208, 210, 212, 213, 207, 207, 212, 211, 215, 212, 215, 214, 215, 214, 217, 218, 216, 218, 216, 215, 215, 217, 215, 214, 217, 220, 220, 219, 217, 220, 219, 219, 217, 219, 220, 220, 221, 220, 217, 220, 218, 222, 220, 220, 219, 221, 217, 221, 219, 216, 221, 220, 221, 220, 221, 221, 220, 219, 220, 220, 222, 221, 223, 224, 225, 223, 220, 219, 221, 225, 224, 224, 223, 223, 225, 225, 224, 222, 221, 220, 222, 221, 222, 224, 221, 226, 224, 223, 219, 219, 220, 220, 220, 221, 220, 220, 223, 221, 221, 217, 220, 222, 223, 221, 220, 223, 224, 224, 224, 224, 224, 224, 223, 224, 223, 224, 222, 223, 223, 225, 222, 221, 224, 220, 222, 225, 224, 223, 221, 223, 226, 222, 223, 222, 222, 221, 224, 223, 222, 223, 223, 222, 223, 221, 221, 219, 224, 221, 222, 220, 220, 222, 221, 221, 221, 223, 222, 223, 219, 220, 219, 218, 220, 220, 222, 224, 221, 221, 222, 223, 223, 222, 218, 223, 220, 216, 219, 219, 218, 222, 223, 219, 221, 222, 224, 224, 224, 221, 220, 220, 222, 222, 224, 221, 221, 219, 222, 221, 223, 221, 220, 220, 225, 219, 222, 221, 220, 222, 220, 218, 218, 217, 215, 222, 215, 216, 217, 215, 220, 220, 222, 217, 214, 209, 193, 204, 204, 197, 203, 102, 192, 201, 202, 203, 201, 201, 201, 204, 205, 205, 206, 206, 207, 206, 203, 209, 205, 208, 207, 211, 210, 209, 208, 207, 212, 209, 209, 213, 210, 212, 212, 210, 212, 212, 214, 213, 216, 216, 213, 214, 215, 216, 217, 220, 217, 215, 218, 213, 215, 215, 218, 220, 221, 220, 217, 222, 221, 220, 220, 221, 220, 219, 221, 221, 219, 221, 219, 221, 221, 217, 216, 219, 220, 222, 219, 219, 220, 221, 222, 219, 222, 222, 221, 220, 221, 221, 221, 223, 225, 225, 223, 221, 220, 220, 222, 225, 225, 224, 224, 221, 225, 225, 226, 223, 222, 223, 224, 224, 222, 224, 225, 225, 227, 223, 223, 222, 220, 221, 222, 222, 221, 218, 222, 220, 218, 220, 221, 222, 222, 221, 222, 222, 224, 224, 225, 223, 221, 223, 222, 225, 224, 224, 223, 223, 224, 221, 221, 219, 223, 223, 225, 226, 225, 223, 222, 225, 224, 223, 223, 223, 225, 226, 225, 223, 225, 221, 223, 223, 223, 221, 221, 220, 224, 223, 220, 221, 220, 223, 223, 221, 222, 221, 223, 223, 221, 221, 220, 223, 221, 221, 222, 221, 221, 220, 222, 223, 224, 219, 221, 223, 221, 217, 222, 222, 221, 225, 223, 222, 221, 223, 223, 223, 224, 223, 223, 220, 220, 223, 222, 220, 223, 223, 222, 222, 219, 221, 221, 221, 225, 223, 222, 220, 220, 222, 218, 220, 218, 217, 214, 220, 218, 216, 217, 218, 220, 218, 218, 218, 212, 205, 186, 208, 203, 198, 201, 89, 191, 204, 202, 202, 200, 203, 203, 204, 203, 205, 203, 205, 206, 205, 203, 205, 207, 208, 207, 212, 208, 210, 210, 209, 209, 207, 211, 212, 213, 208, 212, 213, 212, 210, 213, 216, 217, 211, 213, 214, 216, 217, 215, 218, 219, 219, 218, 217, 218, 214, 217, 220, 221, 223, 217, 219, 221, 222, 221, 223, 219, 220, 222, 222, 221, 219, 220, 224, 221, 221, 218, 220, 222, 222, 222, 220, 218, 219, 220, 218, 223, 223, 220, 219, 221, 223, 222, 223, 223, 223, 225, 219, 220, 219, 223, 222, 222, 224, 225, 224, 225, 225, 226, 223, 221, 223, 223, 225, 223, 223, 225, 226, 224, 225, 221, 222, 222, 221, 223, 220, 221, 220, 222, 222, 223, 222, 221, 223, 222, 224, 225, 222, 221, 224, 225, 224, 223, 223, 221, 222, 224, 223, 223, 224, 222, 224, 223, 223, 224, 225, 226, 225, 224, 224, 223, 226, 225, 225, 223, 225, 226, 227, 224, 226, 224, 225, 224, 221, 223, 222, 222, 222, 223, 222, 222, 221, 222, 221, 225, 222, 222, 221, 222, 224, 223, 223, 219, 222, 224, 220, 223, 223, 223, 220, 224, 222, 222, 222, 222, 224, 222, 224, 220, 220, 225, 224, 223, 223, 222, 221, 224, 223, 224, 222, 221, 221, 223, 221, 223, 221, 220, 222, 222, 221, 219, 219, 221, 218, 223, 224, 222, 221, 223, 222, 221, 218, 218, 216, 217, 219, 215, 217, 219, 220, 222, 219, 225, 219, 214, 208, 185, 206, 205, 201, 200, 94, 193, 203, 204, 204, 203, 205, 202, 203, 205, 207, 204, 207, 207, 204, 207, 204, 210, 207, 208, 209, 207, 207, 206, 208, 208, 213, 212, 209, 212, 212, 211, 214, 211, 212, 214, 214, 215, 216, 215, 214, 218, 218, 216, 219, 218, 218, 217, 219, 217, 217, 218, 221, 219, 219, 220, 220, 221, 220, 220, 222, 219, 223, 221, 223, 223, 222, 221, 223, 220, 220, 218, 221, 222, 222, 221, 221, 220, 219, 220, 218, 221, 223, 224, 222, 220, 224, 224, 224, 222, 222, 227, 220, 220, 221, 223, 225, 225, 224, 225, 224, 226, 224, 224, 225, 223, 224, 223, 222, 224, 222, 224, 222, 223, 222, 222, 223, 224, 226, 223, 224, 223, 222, 221, 224, 225, 221, 224, 224, 222, 225, 224, 223, 223, 225, 226, 223, 223, 222, 223, 221, 222, 224, 224, 224, 224, 226, 226, 225, 225, 226, 226, 227, 226, 223, 224, 225, 225, 224, 226, 225, 225, 227, 226, 225, 225, 222, 222, 224, 225, 224, 222, 221, 221, 220, 222, 222, 225, 224, 223, 224, 221, 222, 223, 225, 224, 222, 222, 224, 225, 223, 224, 222, 222, 223, 224, 224, 224, 222, 222, 224, 222, 222, 223, 220, 223, 221, 223, 223, 222, 224, 224, 224, 226, 224, 222, 220, 223, 220, 225, 222, 221, 223, 222, 224, 223, 222, 219, 220, 222, 226, 222, 224, 224, 219, 221, 221, 220, 216, 218, 217, 218, 217, 219, 222, 220, 222, 223, 220, 215, 207, 190, 203, 198, 196, 200, 97, 199, 205, 207, 205, 203, 206, 205, 205, 204, 206, 204, 207, 205, 210, 211, 208, 211, 210, 212, 211, 203, 209, 204, 207, 207, 209, 209, 207, 213, 211, 214, 213, 212, 209, 214, 215, 219, 216, 214, 216, 217, 218, 221, 220, 218, 219, 215, 218, 216, 217, 217, 221, 222, 223, 222, 220, 222, 220, 222, 222, 221, 223, 222, 222, 220, 220, 220, 223, 220, 219, 220, 220, 221, 218, 222, 219, 220, 220, 224, 224, 224, 224, 223, 222, 222, 226, 224, 223, 224, 224, 225, 224, 219, 221, 223, 226, 222, 225, 224, 224, 225, 226, 225, 223, 224, 223, 224, 222, 224, 224, 224, 223, 223, 222, 224, 224, 220, 225, 224, 224, 222, 224, 222, 225, 225, 224, 225, 224, 223, 225, 223, 223, 225, 227, 227, 223, 225, 221, 225, 223, 223, 223, 224, 226, 226, 226, 227, 226, 226, 226, 227, 228, 226, 223, 224, 225, 227, 225, 227, 227, 225, 227, 225, 224, 223, 222, 225, 226, 224, 223, 224, 222, 224, 222, 222, 224, 224, 225, 223, 224, 222, 220, 224, 224, 224, 224, 220, 224, 224, 226, 222, 223, 224, 222, 225, 223, 224, 223, 222, 225, 225, 223, 223, 225, 222, 224, 224, 223, 224, 225, 224, 225, 224, 226, 219, 221, 222, 222, 224, 224, 220, 223, 222, 223, 224, 224, 219, 224, 224, 225, 224, 223, 222, 224, 221, 220, 221, 217, 220, 216, 216, 221, 217, 221, 218, 224, 220, 218, 216, 209, 194, 202, 203, 200, 203, 93, 199, 205, 201, 206, 206, 207, 205, 207, 209, 208, 206, 210, 208, 210, 212, 210, 210, 210, 209, 213, 209, 208, 210, 208, 208, 208, 209, 211, 212, 213, 212, 212, 214, 211, 216, 217, 218, 216, 218, 216, 218, 217, 218, 219, 216, 221, 216, 219, 218, 219, 220, 220, 221, 223, 222, 222, 221, 224, 224, 222, 222, 224, 224, 224, 223, 220, 222, 222, 223, 219, 220, 218, 217, 219, 222, 219, 218, 222, 222, 225, 224, 223, 221, 224, 224, 224, 224, 225, 224, 224, 224, 222, 220, 221, 223, 223, 225, 223, 226, 224, 224, 225, 224, 224, 224, 225, 224, 225, 224, 225, 223, 223, 225, 225, 223, 222, 224, 224, 223, 224, 222, 223, 223, 224, 224, 224, 224, 225, 226, 226, 224, 224, 226, 227, 226, 225, 225, 224, 223, 225, 223, 224, 224, 224, 226, 226, 226, 227, 226, 226, 227, 225, 225, 224, 225, 227, 227, 228, 225, 225, 223, 226, 226, 224, 224, 222, 223, 225, 225, 224, 221, 222, 223, 223, 223, 224, 225, 225, 224, 225, 223, 223, 224, 225, 224, 223, 224, 224, 224, 227, 225, 223, 224, 223, 224, 225, 223, 224, 224, 223, 225, 223, 222, 221, 223, 222, 222, 222, 223, 223, 222, 226, 224, 224, 221, 222, 222, 223, 226, 221, 222, 223, 224, 224, 223, 222, 217, 219, 223, 224, 225, 223, 224, 222, 223, 219, 219, 220, 217, 219, 215, 217, 215, 220, 220, 223, 220, 220, 218, 210, 193, 203, 203, 201, 202, 100, 198, 207, 202, 202, 206, 207, 204, 207, 211, 207, 210, 211, 211, 210, 212, 213, 209, 212, 211, 212, 212, 210, 210, 212, 210, 209, 210, 210, 212, 210, 215, 213, 213, 217, 217, 218, 217, 215, 218, 217, 218, 223, 220, 217, 216, 220, 215, 220, 220, 220, 222, 222, 220, 221, 221, 218, 223, 223, 223, 223, 224, 223, 222, 223, 222, 221, 222, 221, 222, 217, 220, 220, 219, 222, 222, 218, 219, 222, 224, 224, 223, 220, 224, 222, 225, 225, 225, 224, 223, 225, 223, 225, 220, 221, 224, 225, 224, 224, 225, 223, 225, 224, 227, 224, 224, 226, 227, 227, 225, 224, 224, 221, 224, 225, 224, 222, 224, 225, 226, 224, 224, 225, 222, 225, 225, 224, 223, 224, 225, 226, 224, 225, 227, 229, 228, 229, 225, 224, 223, 222, 224, 223, 223, 223, 224, 225, 227, 227, 225, 226, 226, 229, 227, 226, 224, 226, 224, 225, 226, 225, 227, 228, 228, 225, 224, 224, 225, 224, 224, 225, 223, 224, 226, 224, 225, 225, 224, 225, 226, 227, 223, 222, 225, 225, 224, 224, 222, 222, 223, 226, 224, 222, 223, 224, 223, 225, 226, 224, 224, 224, 223, 224, 220, 220, 219, 224, 223, 224, 224, 225, 224, 224, 223, 224, 223, 221, 222, 218, 224, 220, 223, 223, 223, 224, 225, 222, 220, 221, 224, 224, 225, 224, 223, 224, 222, 222, 219, 217, 219, 220, 216, 222, 220, 221, 220, 219, 222, 219, 214, 208, 193, 204, 203, 204, 204, 102, 200, 203, 202, 203, 207, 209, 207, 210, 208, 211, 208, 208, 210, 210, 211, 215, 208, 215, 213, 216, 212, 209, 212, 210, 211, 210, 210, 210, 214, 212, 215, 211, 213, 218, 216, 219, 218, 218, 216, 216, 220, 221, 220, 217, 218, 216, 217, 215, 221, 218, 222, 220, 225, 224, 221, 222, 224, 223, 223, 221, 223, 223, 222, 223, 221, 220, 219, 221, 222, 217, 219, 219, 220, 222, 219, 221, 221, 220, 221, 223, 225, 223, 224, 225, 228, 225, 225, 224, 225, 227, 225, 226, 222, 223, 224, 226, 223, 225, 227, 227, 225, 226, 226, 222, 224, 227, 226, 226, 226, 223, 223, 223, 224, 225, 224, 224, 224, 223, 226, 224, 225, 224, 225, 224, 227, 222, 223, 224, 224, 225, 225, 226, 225, 228, 228, 228, 227, 226, 224, 227, 224, 226, 225, 226, 225, 227, 228, 227, 225, 226, 229, 228, 227, 224, 225, 227, 224, 227, 226, 227, 226, 227, 229, 226, 224, 226, 222, 226, 226, 223, 223, 224, 225, 224, 227, 225, 223, 227, 226, 227, 223, 222, 223, 224, 225, 223, 224, 222, 223, 226, 226, 224, 225, 223, 225, 224, 225, 224, 223, 226, 225, 224, 221, 223, 220, 224, 224, 227, 224, 223, 224, 224, 224, 222, 225, 223, 225, 226, 223, 222, 224, 225, 223, 223, 224, 222, 220, 224, 225, 224, 225, 223, 223, 224, 222, 222, 220, 220, 219, 220, 221, 219, 223, 221, 222, 221, 222, 217, 217, 208, 194, 205, 201, 202, 203, 102, 198, 205, 202, 201, 206, 206, 208, 212, 208, 210, 205, 206, 210, 211, 214, 213, 213, 214, 211, 212, 213, 211, 210, 213, 214, 211, 214, 212, 212, 213, 212, 214, 215, 219, 217, 218, 219, 217, 217, 219, 219, 219, 219, 220, 219, 220, 220, 218, 219, 218, 222, 222, 223, 223, 222, 224, 221, 224, 221, 222, 224, 221, 224, 223, 221, 221, 220, 220, 220, 218, 219, 220, 222, 221, 219, 222, 222, 222, 222, 225, 224, 224, 223, 224, 225, 224, 225, 226, 224, 226, 225, 224, 225, 225, 226, 226, 226, 226, 227, 226, 225, 226, 226, 224, 224, 224, 226, 225, 224, 225, 223, 226, 226, 226, 224, 224, 226, 226, 226, 226, 223, 224, 226, 224, 225, 224, 224, 225, 224, 226, 225, 225, 226, 228, 229, 229, 225, 227, 226, 226, 226, 227, 227, 225, 226, 228, 226, 226, 224, 225, 229, 227, 226, 221, 223, 225, 225, 226, 227, 227, 226, 228, 227, 228, 225, 227, 226, 226, 224, 223, 225, 223, 224, 224, 224, 226, 224, 226, 226, 225, 225, 224, 223, 224, 225, 224, 224, 224, 224, 227, 227, 224, 223, 221, 226, 226, 225, 223, 223, 225, 225, 224, 225, 222, 223, 223, 225, 225, 223, 224, 224, 224, 223, 224, 225, 223, 224, 224, 223, 223, 225, 227, 222, 224, 224, 225, 223, 224, 225, 226, 224, 225, 220, 225, 224, 222, 219, 219, 219, 220, 222, 221, 223, 222, 222, 221, 222, 220, 213, 208, 195, 207, 200, 201, 202, 99, 197, 203, 202, 204, 206, 204, 207, 211, 214, 212, 209, 206, 207, 213, 213, 215, 214, 215, 216, 212, 214, 215, 214, 213, 214, 211, 212, 213, 214, 216, 213, 213, 216, 217, 219, 220, 216, 218, 216, 218, 218, 221, 220, 221, 220, 221, 221, 220, 221, 222, 223, 223, 224, 222, 220, 224, 224, 224, 222, 223, 223, 221, 224, 223, 223, 223, 221, 223, 220, 220, 219, 219, 222, 223, 222, 223, 220, 221, 226, 224, 224, 224, 223, 226, 227, 226, 226, 226, 226, 227, 227, 224, 226, 225, 227, 226, 226, 226, 228, 226, 226, 227, 225, 226, 224, 224, 226, 225, 224, 224, 225, 226, 227, 227, 225, 224, 226, 224, 225, 225, 225, 225, 225, 225, 225, 225, 226, 226, 224, 224, 227, 225, 228, 229, 229, 228, 227, 227, 228, 226, 227, 227, 225, 225, 225, 226, 224, 225, 224, 225, 228, 229, 227, 224, 222, 226, 223, 227, 225, 225, 227, 227, 228, 228, 226, 226, 226, 227, 225, 221, 225, 222, 222, 225, 224, 224, 224, 225, 226, 227, 225, 224, 224, 223, 224, 224, 223, 224, 222, 226, 226, 226, 221, 221, 227, 226, 224, 224, 223, 225, 224, 227, 224, 219, 224, 226, 225, 225, 222, 222, 225, 223, 222, 225, 224, 225, 222, 224, 216, 220, 223, 223, 222, 226, 225, 224, 222, 225, 224, 224, 220, 221, 221, 224, 224, 221, 224, 221, 222, 221, 222, 221, 221, 219, 223, 220, 219, 217, 212, 205, 195, 207, 204, 202, 201, 105, 198, 204, 202, 203, 205, 207, 209, 210, 213, 211, 205, 208, 212, 212, 211, 215, 216, 213, 214, 211, 212, 213, 215, 214, 214, 211, 213, 213, 216, 215, 216, 215, 217, 217, 218, 220, 220, 220, 220, 220, 219, 219, 221, 222, 220, 221, 223, 221, 219, 223, 224, 222, 221, 223, 221, 221, 224, 222, 223, 224, 223, 223, 226, 225, 223, 223, 224, 224, 224, 219, 221, 219, 222, 223, 224, 222, 223, 222, 226, 226, 226, 223, 225, 226, 226, 227, 225, 225, 225, 227, 226, 223, 225, 224, 226, 225, 224, 225, 227, 226, 227, 227, 225, 225, 226, 227, 226, 226, 224, 225, 226, 226, 226, 226, 225, 223, 225, 227, 225, 226, 224, 226, 227, 226, 227, 226, 227, 227, 228, 226, 226, 227, 226, 228, 229, 229, 228, 226, 228, 227, 229, 228, 226, 224, 226, 227, 227, 227, 228, 228, 228, 228, 227, 226, 224, 225, 226, 226, 227, 225, 227, 227, 228, 229, 227, 226, 225, 227, 225, 224, 222, 222, 225, 224, 225, 224, 224, 227, 227, 226, 225, 224, 224, 225, 226, 223, 223, 224, 225, 228, 227, 225, 223, 224, 225, 226, 223, 222, 224, 223, 226, 226, 223, 224, 222, 223, 226, 224, 223, 223, 224, 225, 225, 224, 224, 224, 225, 227, 221, 219, 225, 224, 225, 225, 225, 224, 224, 227, 225, 224, 220, 223, 222, 222, 225, 223, 219, 222, 220, 222, 222, 220, 220, 223, 222, 221, 222, 220, 214, 205, 198, 203, 207, 201, 205, 92, 196, 203, 205, 204, 204, 212, 212, 211, 213, 208, 203, 207, 212, 213, 214, 216, 216, 213, 212, 214, 214, 213, 216, 214, 214, 213, 212, 213, 217, 214, 216, 214, 218, 219, 217, 219, 220, 222, 220, 219, 218, 220, 220, 223, 219, 222, 221, 220, 221, 222, 224, 224, 224, 221, 222, 222, 222, 222, 223, 223, 222, 224, 226, 225, 225, 224, 225, 224, 224, 222, 218, 221, 224, 223, 223, 225, 222, 225, 226, 227, 226, 224, 225, 226, 226, 226, 226, 225, 227, 227, 225, 226, 225, 226, 225, 224, 227, 226, 227, 226, 226, 227, 227, 225, 226, 227, 225, 225, 226, 226, 226, 227, 227, 227, 225, 224, 224, 228, 225, 226, 226, 225, 226, 227, 227, 225, 228, 228, 228, 226, 227, 227, 226, 227, 228, 227, 228, 228, 228, 228, 228, 226, 227, 224, 229, 227, 227, 225, 226, 227, 227, 230, 228, 226, 226, 226, 224, 227, 226, 224, 226, 226, 229, 228, 227, 227, 226, 225, 227, 223, 223, 223, 225, 226, 226, 226, 226, 227, 227, 225, 226, 225, 224, 226, 225, 223, 224, 223, 225, 225, 227, 223, 224, 225, 225, 225, 227, 224, 224, 222, 227, 225, 225, 225, 225, 226, 225, 225, 224, 222, 223, 225, 224, 225, 225, 225, 227, 227, 221, 223, 224, 227, 227, 226, 225, 225, 224, 225, 225, 225, 223, 222, 221, 224, 225, 223, 220, 220, 223, 220, 221, 221, 220, 224, 221, 224, 220, 218, 213, 207, 199, 204, 202, 203, 209, 120, 201, 206, 204, 205, 205, 209, 211, 212, 212, 210, 206, 208, 209, 214, 215, 212, 212, 211, 211, 215, 214, 216, 215, 214, 214, 214, 213, 216, 218, 215, 213, 216, 218, 219, 222, 218, 222, 220, 222, 221, 221, 219, 222, 224, 219, 223, 222, 221, 219, 221, 221, 226, 224, 223, 220, 222, 221, 223, 222, 224, 221, 223, 225, 225, 225, 224, 224, 225, 224, 223, 223, 221, 224, 223, 222, 222, 222, 225, 225, 226, 226, 224, 223, 225, 227, 225, 224, 224, 226, 227, 226, 226, 223, 227, 227, 226, 227, 227, 226, 226, 227, 226, 226, 224, 225, 226, 225, 226, 224, 225, 224, 225, 226, 227, 226, 226, 227, 227, 225, 226, 225, 225, 226, 229, 227, 226, 227, 226, 227, 226, 226, 226, 227, 226, 230, 229, 227, 228, 228, 229, 229, 227, 226, 225, 227, 226, 228, 226, 225, 229, 229, 227, 228, 226, 226, 229, 227, 227, 225, 227, 227, 228, 229, 228, 228, 228, 228, 226, 227, 224, 221, 223, 225, 225, 225, 226, 227, 228, 226, 227, 227, 225, 224, 227, 226, 225, 223, 223, 223, 226, 226, 226, 222, 225, 227, 224, 227, 225, 224, 224, 226, 226, 224, 226, 224, 228, 225, 222, 221, 222, 221, 226, 226, 224, 225, 227, 226, 227, 225, 225, 223, 226, 227, 225, 226, 223, 224, 226, 226, 225, 224, 224, 224, 224, 224, 223, 222, 222, 220, 219, 220, 223, 221, 222, 222, 222, 220, 220, 217, 208, 201, 204, 204, 202, 208, 124, 208, 201, 204, 210, 207, 211, 207, 215, 215, 214, 210, 208, 210, 212, 213, 211, 212, 212, 209, 216, 214, 214, 212, 214, 216, 214, 211, 216, 215, 212, 216, 218, 218, 218, 221, 221, 219, 220, 221, 222, 222, 219, 221, 224, 221, 224, 222, 224, 221, 221, 222, 224, 221, 221, 222, 219, 222, 223, 224, 224, 221, 223, 224, 224, 225, 224, 224, 222, 222, 223, 224, 221, 223, 222, 225, 223, 225, 225, 226, 225, 226, 225, 224, 227, 226, 224, 223, 225, 226, 226, 227, 227, 226, 227, 226, 227, 227, 227, 226, 227, 227, 227, 228, 226, 225, 227, 227, 227, 225, 225, 222, 226, 227, 227, 225, 226, 227, 226, 227, 226, 224, 225, 227, 227, 227, 224, 226, 226, 225, 227, 227, 227, 226, 228, 227, 228, 228, 227, 228, 229, 228, 228, 227, 225, 227, 228, 225, 226, 226, 227, 229, 227, 228, 228, 228, 228, 227, 228, 227, 226, 228, 227, 227, 228, 228, 227, 225, 225, 228, 225, 223, 224, 225, 224, 225, 225, 226, 226, 225, 224, 226, 225, 222, 226, 227, 225, 224, 220, 223, 223, 224, 227, 225, 226, 225, 225, 223, 223, 222, 225, 224, 225, 226, 226, 225, 225, 224, 221, 223, 222, 223, 226, 227, 224, 224, 226, 226, 227, 226, 226, 224, 228, 227, 227, 227, 225, 224, 226, 226, 227, 226, 225, 227, 225, 226, 221, 220, 220, 223, 222, 220, 221, 221, 221, 222, 222, 223, 219, 217, 209, 204, 207, 205, 202, 209, 135, 204, 203, 207, 208, 212, 210, 212, 214, 215, 213, 209, 209, 212, 212, 213, 212, 210, 211, 210, 213, 213, 213, 215, 215, 216, 213, 214, 213, 217, 214, 217, 217, 215, 216, 222, 222, 221, 220, 219, 223, 221, 221, 223, 223, 224, 224, 224, 223, 221, 221, 223, 225, 219, 224, 223, 222, 225, 222, 222, 223, 222, 224, 225, 225, 225, 225, 223, 226, 223, 222, 223, 224, 224, 226, 225, 223, 224, 225, 227, 225, 226, 225, 225, 225, 226, 225, 221, 225, 225, 224, 227, 225, 227, 227, 227, 227, 228, 227, 226, 225, 227, 227, 228, 227, 225, 226, 227, 227, 223, 225, 223, 226, 227, 226, 225, 226, 227, 225, 227, 226, 226, 226, 228, 228, 228, 226, 226, 226, 228, 226, 226, 227, 227, 229, 228, 228, 228, 227, 227, 228, 229, 228, 227, 227, 229, 227, 223, 225, 226, 227, 226, 229, 228, 227, 227, 227, 227, 228, 226, 228, 228, 228, 228, 228, 228, 227, 226, 228, 227, 225, 225, 222, 224, 224, 227, 225, 226, 226, 226, 227, 223, 225, 226, 225, 226, 226, 224, 224, 224, 222, 226, 227, 226, 226, 224, 225, 225, 223, 224, 224, 223, 224, 223, 224, 224, 226, 226, 224, 225, 223, 225, 225, 227, 225, 225, 226, 225, 228, 227, 225, 226, 227, 228, 228, 227, 225, 224, 226, 224, 225, 225, 225, 228, 226, 226, 224, 223, 222, 221, 222, 224, 221, 222, 222, 221, 222, 219, 217, 214, 211, 206, 208, 200, 204, 210, 120, 202, 207, 208, 208, 210, 208, 210, 209, 212, 212, 211, 211, 212, 214, 213, 208, 211, 214, 213, 213, 211, 213, 215, 210, 212, 215, 217, 214, 218, 217, 221, 218, 217, 218, 225, 221, 222, 222, 219, 223, 223, 224, 224, 225, 225, 225, 226, 224, 224, 223, 225, 225, 221, 224, 223, 224, 224, 226, 224, 224, 222, 224, 224, 224, 226, 226, 223, 224, 224, 224, 224, 225, 226, 225, 226, 225, 224, 225, 225, 225, 225, 224, 225, 226, 226, 225, 225, 224, 225, 225, 224, 226, 226, 225, 226, 227, 228, 225, 226, 227, 227, 227, 228, 227, 226, 228, 229, 227, 226, 225, 225, 228, 226, 226, 226, 227, 228, 225, 226, 227, 226, 227, 227, 228, 228, 228, 228, 228, 230, 226, 227, 227, 228, 228, 228, 228, 228, 228, 227, 228, 228, 228, 228, 228, 228, 228, 225, 224, 225, 225, 228, 229, 228, 228, 228, 228, 230, 230, 228, 227, 226, 227, 229, 229, 225, 227, 228, 224, 226, 227, 223, 225, 226, 225, 225, 224, 224, 224, 226, 227, 224, 225, 224, 225, 227, 227, 225, 223, 222, 224, 225, 225, 223, 224, 225, 226, 225, 224, 223, 224, 226, 225, 222, 224, 225, 227, 228, 226, 224, 224, 224, 227, 226, 225, 225, 227, 224, 228, 226, 225, 227, 226, 228, 227, 226, 224, 226, 225, 226, 225, 225, 225, 225, 224, 227, 225, 223, 223, 219, 221, 221, 222, 221, 223, 220, 218, 218, 215, 219, 212, 205, 207, 202, 201, 206, 112, 204, 205, 211, 207, 211, 208, 210, 208, 211, 212, 213, 212, 211, 214, 214, 212, 213, 215, 210, 212, 211, 212, 212, 213, 217, 215, 216, 213, 217, 220, 220, 219, 215, 217, 223, 224, 221, 222, 222, 224, 226, 224, 224, 224, 225, 223, 227, 225, 223, 224, 226, 224, 223, 222, 224, 227, 225, 226, 225, 224, 224, 226, 225, 223, 227, 224, 224, 224, 224, 222, 224, 224, 224, 225, 227, 225, 226, 227, 228, 226, 225, 225, 225, 226, 226, 225, 226, 224, 225, 226, 226, 226, 228, 226, 228, 227, 229, 227, 226, 227, 227, 227, 227, 227, 226, 225, 229, 227, 226, 227, 226, 229, 227, 227, 226, 228, 227, 229, 226, 226, 227, 226, 228, 227, 228, 227, 228, 228, 230, 228, 228, 225, 227, 228, 229, 229, 229, 228, 228, 228, 227, 229, 228, 228, 229, 228, 227, 226, 225, 228, 229, 229, 228, 228, 227, 228, 230, 229, 229, 225, 226, 225, 228, 228, 225, 226, 227, 226, 225, 226, 225, 224, 226, 227, 225, 223, 225, 226, 224, 225, 221, 224, 225, 224, 226, 223, 224, 223, 225, 226, 225, 225, 224, 225, 226, 226, 225, 222, 224, 223, 226, 224, 225, 225, 225, 227, 228, 227, 226, 224, 227, 227, 227, 226, 225, 226, 226, 226, 227, 225, 228, 227, 226, 226, 226, 226, 223, 224, 226, 225, 224, 225, 226, 225, 225, 220, 222, 221, 222, 220, 221, 222, 221, 221, 220, 220, 221, 219, 217, 211, 205, 209, 203, 204, 206, 113, 202, 211, 209, 210, 207, 207, 209, 208, 215, 214, 214, 212, 213, 215, 212, 213, 214, 216, 212, 212, 216, 215, 213, 216, 220, 215, 217, 216, 218, 222, 219, 220, 216, 217, 224, 222, 220, 220, 221, 225, 226, 223, 223, 224, 224, 225, 224, 225, 224, 225, 224, 226, 225, 225, 226, 225, 226, 225, 225, 223, 225, 226, 226, 226, 227, 224, 225, 226, 226, 224, 226, 226, 224, 225, 226, 224, 226, 226, 227, 227, 225, 226, 226, 226, 227, 226, 224, 224, 225, 228, 229, 226, 227, 226, 228, 227, 227, 227, 226, 228, 227, 228, 228, 227, 227, 226, 229, 227, 227, 227, 226, 228, 230, 228, 226, 227, 227, 227, 227, 226, 227, 228, 227, 227, 229, 227, 228, 228, 230, 229, 228, 227, 227, 228, 228, 228, 227, 227, 227, 228, 227, 230, 228, 228, 229, 228, 229, 227, 226, 227, 229, 229, 227, 228, 228, 228, 230, 229, 227, 227, 225, 225, 227, 226, 222, 225, 226, 226, 226, 226, 224, 223, 225, 226, 227, 224, 225, 225, 224, 221, 221, 222, 225, 225, 224, 225, 224, 226, 224, 226, 226, 226, 226, 226, 227, 227, 228, 225, 225, 226, 228, 227, 226, 227, 224, 227, 227, 226, 223, 226, 226, 226, 226, 224, 225, 225, 227, 227, 229, 228, 227, 226, 228, 227, 225, 225, 224, 225, 226, 225, 225, 225, 227, 226, 223, 223, 225, 220, 222, 222, 223, 222, 222, 221, 220, 222, 219, 219, 218, 209, 205, 206, 202, 201, 204, 109, 204, 208, 213, 210, 203, 206, 212, 208, 214, 214, 211, 212, 214, 215, 213, 216, 215, 213, 214, 213, 217, 216, 218, 216, 220, 216, 217, 218, 220, 224, 221, 219, 214, 218, 222, 220, 222, 219, 221, 223, 225, 222, 221, 224, 224, 224, 225, 227, 226, 224, 225, 226, 225, 225, 224, 225, 225, 225, 225, 225, 226, 226, 228, 227, 225, 225, 225, 225, 226, 225, 226, 225, 226, 226, 227, 224, 226, 226, 227, 228, 226, 226, 224, 225, 225, 225, 225, 224, 225, 227, 227, 225, 227, 227, 226, 228, 229, 227, 227, 227, 227, 229, 227, 227, 227, 227, 228, 229, 228, 228, 228, 229, 229, 227, 226, 228, 227, 229, 228, 227, 228, 228, 229, 228, 228, 228, 227, 229, 229, 230, 229, 226, 227, 229, 229, 228, 227, 228, 228, 229, 229, 228, 227, 227, 229, 229, 228, 228, 227, 228, 230, 229, 228, 226, 226, 229, 230, 227, 226, 226, 226, 226, 227, 226, 223, 225, 227, 227, 225, 226, 224, 221, 224, 225, 228, 225, 226, 225, 224, 222, 222, 220, 225, 223, 224, 223, 222, 226, 225, 227, 227, 228, 226, 225, 228, 226, 226, 227, 226, 226, 227, 228, 226, 225, 226, 228, 227, 224, 223, 227, 227, 226, 225, 223, 224, 225, 227, 228, 230, 228, 227, 228, 228, 227, 228, 225, 224, 226, 225, 226, 226, 225, 223, 224, 225, 222, 224, 221, 224, 222, 224, 222, 222, 224, 221, 219, 219, 220, 218, 210, 211, 209, 206, 201, 205, 101, 204, 209, 211, 210, 204, 207, 210, 208, 211, 214, 211, 210, 216, 215, 213, 216, 216, 217, 215, 217, 217, 216, 216, 217, 221, 219, 217, 217, 220, 222, 220, 218, 214, 215, 222, 218, 220, 221, 221, 220, 223, 222, 224, 225, 224, 225, 226, 225, 226, 224, 227, 225, 225, 223, 224, 224, 225, 223, 225, 224, 226, 226, 227, 226, 225, 225, 225, 224, 226, 225, 226, 225, 226, 227, 226, 225, 226, 225, 228, 227, 227, 224, 225, 224, 224, 224, 225, 226, 226, 228, 228, 227, 227, 226, 227, 227, 227, 228, 225, 226, 227, 228, 228, 228, 227, 228, 229, 228, 228, 228, 227, 227, 229, 228, 227, 227, 227, 227, 228, 228, 227, 228, 228, 228, 228, 227, 229, 230, 230, 229, 227, 228, 227, 228, 227, 228, 229, 229, 229, 230, 228, 228, 228, 227, 229, 228, 229, 227, 228, 228, 229, 230, 228, 226, 226, 229, 228, 229, 226, 226, 225, 227, 227, 227, 224, 225, 225, 227, 227, 228, 225, 224, 223, 226, 226, 227, 226, 226, 225, 223, 222, 222, 223, 223, 221, 224, 222, 223, 224, 227, 227, 227, 227, 227, 227, 229, 227, 225, 226, 225, 227, 225, 224, 226, 226, 227, 228, 227, 225, 226, 226, 226, 226, 225, 225, 226, 228, 228, 228, 227, 227, 228, 227, 228, 228, 228, 227, 227, 226, 226, 224, 225, 225, 224, 222, 223, 222, 224, 226, 224, 222, 224, 222, 226, 223, 222, 220, 221, 217, 209, 208, 207, 202, 199, 206, 96, 203, 213, 211, 209, 206, 208, 209, 214, 214, 211, 215, 215, 213, 213, 210, 218, 218, 217, 218, 215, 216, 215, 217, 218, 221, 220, 218, 220, 223, 221, 218, 216, 216, 215, 218, 220, 221, 220, 222, 221, 223, 221, 224, 223, 224, 226, 227, 225, 227, 225, 225, 226, 227, 225, 226, 224, 223, 225, 225, 226, 225, 226, 225, 225, 227, 224, 223, 224, 226, 227, 227, 226, 226, 227, 228, 225, 226, 226, 227, 227, 227, 226, 226, 226, 225, 225, 226, 225, 227, 228, 227, 228, 226, 227, 228, 228, 229, 228, 227, 227, 228, 229, 228, 228, 226, 227, 228, 229, 228, 228, 228, 229, 229, 227, 227, 227, 227, 229, 227, 228, 226, 228, 228, 229, 229, 229, 229, 229, 230, 230, 228, 226, 228, 227, 228, 228, 228, 229, 228, 230, 230, 229, 228, 229, 230, 229, 230, 229, 229, 229, 229, 228, 228, 227, 227, 229, 229, 228, 227, 225, 226, 228, 229, 225, 226, 225, 227, 228, 228, 226, 224, 224, 225, 226, 227, 228, 228, 226, 226, 224, 223, 224, 223, 220, 223, 221, 221, 221, 225, 227, 227, 226, 227, 226, 229, 228, 228, 226, 226, 227, 229, 226, 227, 225, 225, 227, 227, 226, 224, 226, 227, 226, 227, 226, 225, 226, 229, 230, 228, 228, 227, 227, 229, 228, 227, 226, 226, 228, 227, 224, 225, 225, 224, 224, 226, 224, 224, 224, 226, 227, 225, 224, 224, 224, 223, 221, 218, 220, 218, 212, 209, 210, 204, 202, 205, 107, 204, 211, 213, 213, 208, 210, 211, 214, 212, 213, 213, 214, 216, 213, 215, 214, 217, 216, 214, 212, 213, 216, 214, 215, 220, 222, 221, 218, 224, 223, 219, 216, 216, 217, 218, 218, 220, 219, 221, 221, 222, 222, 222, 224, 226, 226, 226, 225, 227, 225, 227, 225, 226, 225, 227, 223, 224, 225, 225, 227, 227, 226, 224, 225, 225, 225, 222, 224, 226, 226, 226, 225, 226, 227, 227, 227, 226, 226, 228, 226, 228, 225, 225, 226, 226, 226, 226, 225, 226, 227, 226, 227, 227, 226, 226, 228, 228, 227, 227, 228, 229, 229, 229, 227, 228, 228, 228, 228, 228, 228, 228, 229, 229, 226, 227, 227, 228, 229, 228, 227, 227, 229, 229, 230, 229, 228, 228, 228, 229, 229, 228, 227, 227, 228, 229, 227, 228, 228, 228, 229, 229, 229, 228, 229, 230, 230, 230, 228, 228, 229, 229, 228, 228, 228, 229, 229, 230, 227, 226, 226, 226, 227, 228, 225, 227, 227, 228, 228, 228, 226, 223, 224, 226, 226, 226, 227, 227, 225, 225, 226, 223, 223, 225, 224, 223, 222, 221, 221, 225, 225, 228, 226, 227, 227, 229, 228, 228, 226, 226, 227, 227, 225, 224, 225, 223, 227, 228, 227, 226, 224, 227, 227, 227, 228, 228, 227, 229, 228, 229, 227, 227, 227, 228, 229, 226, 223, 225, 225, 226, 225, 226, 223, 225, 226, 227, 225, 223, 224, 224, 226, 223, 226, 225, 224, 221, 222, 220, 219, 217, 215, 212, 211, 203, 207, 208, 114, 202, 211, 210, 211, 209, 207, 211, 215, 217, 215, 217, 218, 218, 216, 215, 214, 218, 219, 214, 216, 210, 212, 214, 216, 218, 220, 220, 218, 223, 221, 220, 222, 220, 220, 222, 222, 223, 221, 219, 221, 221, 223, 221, 224, 226, 226, 227, 225, 226, 226, 225, 225, 225, 225, 226, 225, 224, 226, 227, 227, 225, 226, 224, 226, 224, 223, 224, 225, 225, 225, 225, 224, 226, 226, 227, 227, 227, 228, 228, 227, 226, 225, 225, 225, 225, 225, 225, 226, 227, 228, 228, 227, 227, 225, 225, 227, 227, 227, 226, 227, 228, 228, 228, 227, 227, 229, 228, 228, 226, 228, 228, 228, 230, 228, 227, 228, 228, 229, 229, 228, 228, 227, 230, 230, 229, 228, 228, 229, 228, 228, 227, 226, 227, 229, 228, 228, 229, 228, 229, 229, 230, 228, 229, 229, 229, 229, 230, 228, 227, 227, 229, 229, 229, 228, 230, 230, 231, 229, 227, 226, 225, 227, 229, 226, 227, 227, 228, 227, 226, 225, 224, 225, 226, 228, 228, 226, 226, 227, 227, 227, 222, 224, 225, 226, 227, 223, 223, 223, 225, 223, 227, 227, 227, 227, 228, 227, 229, 226, 226, 227, 227, 227, 226, 226, 226, 228, 228, 227, 226, 227, 228, 229, 228, 227, 227, 226, 228, 228, 229, 227, 227, 225, 227, 228, 227, 225, 226, 228, 227, 226, 225, 221, 225, 226, 227, 226, 224, 222, 225, 225, 226, 227, 225, 224, 222, 220, 220, 221, 218, 212, 212, 212, 208, 210, 210, 125, 204, 213, 210, 211, 211, 210, 209, 214, 216, 215, 215, 214, 217, 218, 215, 218, 217, 217, 216, 216, 214, 216, 214, 218, 220, 222, 218, 220, 222, 221, 219, 221, 220, 221, 221, 222, 222, 219, 221, 222, 223, 224, 222, 224, 225, 226, 228, 225, 226, 226, 228, 226, 227, 226, 226, 224, 225, 227, 227, 225, 225, 226, 226, 225, 223, 223, 225, 224, 225, 225, 226, 226, 226, 227, 227, 227, 227, 228, 228, 227, 228, 227, 226, 227, 227, 228, 226, 227, 227, 228, 228, 228, 228, 226, 226, 226, 227, 227, 225, 227, 226, 228, 228, 228, 227, 229, 228, 228, 225, 227, 227, 229, 230, 229, 228, 226, 228, 229, 229, 228, 228, 228, 230, 229, 230, 228, 229, 228, 230, 228, 228, 228, 228, 230, 230, 230, 229, 228, 229, 231, 229, 229, 229, 230, 228, 230, 230, 229, 227, 227, 229, 228, 229, 230, 230, 230, 231, 229, 227, 227, 226, 227, 229, 226, 222, 218, 212, 207, 203, 199, 200, 205, 212, 218, 221, 223, 226, 226, 224, 226, 221, 225, 225, 225, 227, 226, 224, 224, 225, 223, 224, 226, 226, 225, 227, 228, 228, 226, 225, 229, 228, 229, 227, 227, 225, 228, 228, 228, 227, 228, 226, 227, 227, 228, 228, 227, 228, 230, 228, 227, 226, 226, 228, 227, 227, 225, 227, 228, 227, 227, 225, 222, 226, 226, 227, 226, 225, 225, 225, 227, 228, 226, 227, 222, 222, 223, 223, 221, 218, 214, 215, 211, 210, 209, 212, 117, 204, 213, 211, 210, 210, 209, 210, 214, 215, 211, 214, 215, 218, 217, 215, 217, 217, 221, 219, 219, 214, 217, 217, 218, 218, 219, 220, 221, 221, 220, 220, 222, 221, 222, 223, 223, 222, 223, 222, 225, 225, 226, 225, 224, 224, 228, 228, 227, 227, 227, 228, 225, 226, 225, 226, 226, 226, 227, 228, 225, 226, 227, 227, 223, 221, 224, 226, 225, 225, 226, 226, 226, 227, 228, 228, 227, 227, 227, 228, 228, 228, 227, 228, 228, 228, 228, 226, 229, 227, 228, 227, 229, 228, 227, 227, 227, 226, 227, 226, 228, 227, 230, 228, 227, 227, 228, 229, 228, 226, 226, 228, 229, 229, 229, 229, 227, 228, 228, 230, 229, 229, 228, 230, 228, 230, 230, 228, 229, 231, 229, 228, 227, 229, 230, 230, 229, 229, 228, 229, 230, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 233, 233, 232, 234, 235, 233, 232, 230, 224, 209, 191, 162, 134, 108, 90, 76, 74, 68, 69, 71, 84, 96, 123, 147, 175, 192, 202, 211, 216, 220, 225, 226, 227, 228, 225, 227, 226, 224, 225, 225, 228, 229, 228, 227, 228, 227, 225, 226, 228, 229, 226, 226, 227, 226, 229, 229, 226, 228, 228, 229, 229, 229, 228, 228, 228, 229, 229, 226, 225, 227, 227, 226, 228, 227, 226, 228, 228, 228, 225, 225, 226, 225, 227, 227, 225, 224, 227, 226, 227, 226, 224, 219, 222, 222, 223, 223, 217, 213, 211, 213, 212, 210, 212, 124, 208, 214, 211, 210, 208, 211, 210, 210, 216, 212, 216, 212, 218, 216, 217, 217, 218, 219, 219, 219, 216, 214, 219, 216, 220, 220, 219, 222, 223, 220, 222, 221, 221, 221, 222, 224, 224, 221, 223, 221, 226, 227, 224, 224, 224, 226, 226, 226, 226, 226, 227, 224, 225, 226, 226, 226, 227, 226, 227, 226, 226, 226, 227, 226, 223, 224, 226, 225, 225, 225, 226, 225, 227, 228, 228, 226, 226, 227, 226, 228, 228, 228, 227, 227, 228, 227, 228, 228, 227, 228, 228, 229, 228, 227, 227, 228, 228, 226, 228, 227, 229, 230, 230, 228, 228, 228, 229, 226, 227, 227, 228, 229, 230, 230, 229, 229, 229, 230, 230, 230, 229, 229, 229, 228, 229, 229, 229, 228, 231, 229, 228, 228, 230, 230, 230, 230, 230, 230, 230, 231, 231, 232, 231, 232, 233, 234, 234, 232, 232, 233, 235, 235, 235, 235, 236, 236, 236, 231, 212, 169, 121, 82, 70, 67, 65, 68, 74, 78, 81, 75, 76, 79, 77, 83, 80, 74, 70, 78, 96, 134, 159, 179, 195, 212, 221, 224, 222, 227, 226, 227, 226, 226, 228, 228, 228, 229, 228, 227, 228, 228, 228, 229, 228, 227, 227, 227, 226, 229, 227, 227, 228, 229, 227, 228, 228, 227, 227, 228, 229, 226, 226, 228, 229, 227, 228, 227, 226, 228, 228, 228, 226, 227, 223, 225, 228, 227, 224, 224, 227, 227, 227, 226, 225, 223, 222, 223, 225, 222, 218, 215, 213, 211, 208, 211, 212, 132, 209, 216, 211, 210, 214, 211, 209, 211, 212, 214, 213, 214, 216, 219, 219, 219, 218, 220, 219, 219, 219, 217, 219, 219, 219, 222, 221, 221, 222, 223, 222, 222, 222, 224, 222, 225, 224, 223, 225, 224, 227, 225, 225, 223, 225, 226, 226, 226, 225, 225, 228, 227, 226, 226, 226, 226, 227, 227, 227, 227, 227, 227, 228, 228, 226, 227, 226, 227, 226, 225, 226, 226, 227, 228, 227, 227, 227, 226, 228, 228, 226, 228, 227, 227, 229, 228, 227, 228, 228, 228, 229, 230, 227, 227, 228, 229, 228, 228, 228, 227, 230, 230, 230, 227, 229, 229, 230, 230, 228, 228, 227, 230, 230, 230, 229, 228, 230, 230, 229, 229, 228, 228, 230, 230, 229, 229, 229, 230, 231, 231, 229, 229, 229, 230, 231, 231, 230, 231, 231, 231, 234, 232, 232, 232, 233, 234, 234, 234, 234, 235, 236, 236, 237, 237, 236, 231, 215, 157, 89, 68, 69, 72, 78, 84, 86, 87, 88, 94, 94, 98, 111, 114, 123, 130, 118, 100, 88, 78, 69, 63, 63, 86, 115, 151, 175, 198, 214, 221, 226, 228, 226, 226, 227, 224, 228, 228, 229, 227, 227, 228, 228, 230, 228, 227, 227, 228, 228, 227, 228, 227, 228, 229, 229, 227, 228, 227, 227, 227, 228, 227, 224, 228, 229, 229, 229, 227, 228, 227, 227, 229, 227, 226, 225, 226, 226, 224, 227, 225, 227, 226, 227, 224, 223, 222, 223, 224, 226, 224, 218, 215, 205, 211, 210, 209, 212, 129, 208, 217, 212, 213, 212, 206, 207, 213, 215, 212, 215, 215, 219, 219, 218, 217, 218, 221, 219, 219, 218, 219, 218, 220, 221, 218, 221, 222, 221, 219, 223, 225, 222, 225, 226, 224, 224, 224, 224, 224, 228, 226, 226, 225, 224, 228, 226, 224, 224, 226, 229, 227, 228, 226, 226, 225, 228, 228, 228, 227, 227, 227, 228, 228, 226, 226, 227, 228, 227, 225, 225, 226, 226, 227, 227, 226, 228, 228, 228, 228, 227, 228, 227, 228, 227, 228, 227, 228, 228, 229, 229, 230, 228, 227, 228, 229, 228, 228, 228, 228, 229, 230, 229, 229, 229, 230, 230, 230, 229, 228, 227, 229, 229, 230, 229, 228, 228, 230, 230, 229, 229, 228, 231, 231, 229, 229, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 231, 232, 232, 232, 232, 232, 231, 232, 233, 233, 233, 233, 234, 234, 235, 236, 235, 232, 227, 203, 117, 73, 75, 96, 129, 147, 132, 103, 92, 102, 120, 146, 164, 181, 188, 200, 206, 210, 208, 207, 193, 168, 138, 93, 81, 73, 65, 72, 97, 127, 160, 198, 215, 226, 227, 227, 226, 226, 229, 229, 228, 227, 226, 227, 227, 230, 228, 227, 227, 227, 228, 229, 229, 229, 229, 228, 230, 229, 226, 226, 229, 229, 229, 226, 226, 227, 229, 228, 228, 229, 227, 227, 228, 226, 226, 224, 225, 227, 227, 226, 226, 222, 227, 225, 226, 225, 223, 224, 225, 226, 226, 224, 217, 213, 209, 210, 211, 209, 214, 124, 209, 216, 215, 215, 213, 215, 210, 216, 217, 217, 212, 217, 218, 220, 218, 218, 219, 219, 219, 219, 218, 222, 220, 219, 220, 216, 220, 221, 223, 222, 224, 224, 224, 226, 228, 226, 225, 224, 226, 227, 227, 227, 226, 224, 224, 226, 226, 224, 226, 226, 228, 226, 226, 226, 224, 224, 228, 229, 228, 227, 228, 227, 228, 227, 227, 225, 227, 229, 228, 226, 226, 225, 227, 224, 225, 225, 228, 227, 229, 228, 228, 227, 227, 228, 229, 228, 227, 226, 228, 229, 229, 229, 227, 228, 228, 229, 229, 229, 228, 228, 230, 230, 230, 230, 229, 230, 229, 228, 228, 228, 228, 230, 230, 230, 229, 229, 228, 229, 229, 229, 229, 229, 230, 231, 230, 229, 228, 230, 231, 231, 231, 230, 230, 231, 231, 231, 231, 230, 231, 232, 231, 231, 229, 230, 230, 232, 232, 233, 233, 232, 235, 234, 231, 224, 205, 110, 74, 86, 156, 201, 192, 146, 101, 105, 145, 178, 201, 215, 222, 226, 226, 224, 228, 229, 230, 230, 230, 228, 222, 209, 177, 125, 85, 77, 63, 78, 94, 116, 164, 206, 225, 226, 227, 226, 226, 229, 229, 228, 228, 228, 226, 227, 227, 227, 227, 228, 229, 229, 227, 228, 229, 229, 229, 229, 227, 227, 229, 229, 229, 228, 226, 228, 229, 229, 229, 228, 227, 227, 229, 227, 228, 224, 226, 227, 226, 228, 225, 224, 225, 224, 225, 224, 224, 224, 225, 226, 224, 223, 218, 213, 216, 211, 209, 210, 215, 141, 211, 216, 213, 217, 212, 212, 212, 215, 216, 218, 213, 217, 219, 217, 217, 219, 220, 219, 220, 222, 219, 220, 218, 219, 220, 217, 220, 222, 222, 223, 225, 224, 225, 227, 227, 226, 225, 222, 225, 227, 226, 226, 224, 224, 224, 225, 226, 226, 227, 226, 226, 229, 229, 227, 225, 226, 226, 228, 227, 227, 227, 227, 227, 228, 226, 227, 227, 228, 228, 227, 225, 226, 225, 228, 227, 226, 227, 227, 228, 229, 228, 228, 227, 228, 229, 229, 228, 227, 228, 229, 230, 230, 227, 228, 228, 229, 229, 229, 229, 229, 229, 230, 230, 229, 228, 230, 230, 230, 228, 228, 229, 230, 229, 230, 229, 228, 229, 230, 230, 228, 229, 229, 229, 230, 230, 229, 229, 229, 231, 231, 230, 230, 228, 230, 232, 231, 229, 230, 231, 232, 233, 230, 230, 230, 231, 232, 231, 232, 232, 233, 234, 232, 226, 213, 147, 82, 95, 182, 217, 204, 155, 104, 122, 176, 210, 223, 226, 230, 230, 230, 230, 228, 228, 228, 230, 229, 229, 232, 232, 231, 228, 217, 187, 125, 81, 71, 72, 89, 100, 139, 194, 218, 224, 226, 228, 229, 229, 228, 229, 225, 225, 225, 228, 228, 227, 228, 230, 230, 228, 228, 229, 230, 230, 229, 227, 228, 229, 229, 229, 227, 228, 227, 229, 229, 228, 229, 226, 227, 228, 228, 226, 226, 227, 227, 227, 225, 225, 225, 224, 223, 225, 226, 222, 225, 227, 225, 223, 223, 218, 212, 213, 213, 210, 210, 215, 128, 210, 215, 218, 218, 214, 208, 213, 215, 214, 212, 216, 215, 219, 218, 215, 218, 218, 224, 223, 223, 220, 218, 217, 222, 216, 219, 223, 224, 224, 225, 224, 223, 224, 224, 225, 227, 224, 224, 224, 226, 227, 226, 226, 224, 224, 226, 223, 225, 225, 225, 226, 229, 228, 228, 226, 226, 228, 228, 228, 228, 227, 228, 228, 228, 228, 226, 228, 228, 228, 228, 226, 226, 227, 227, 228, 226, 226, 227, 229, 229, 229, 227, 227, 227, 228, 228, 228, 228, 227, 229, 229, 229, 228, 228, 228, 229, 230, 229, 228, 228, 230, 230, 230, 229, 228, 230, 231, 230, 229, 229, 229, 230, 230, 230, 229, 229, 229, 229, 230, 229, 229, 228, 227, 228, 230, 229, 229, 230, 231, 232, 230, 229, 228, 231, 231, 231, 231, 230, 231, 232, 233, 232, 231, 231, 231, 231, 232, 232, 233, 233, 232, 228, 217, 191, 76, 83, 181, 220, 212, 167, 103, 119, 185, 222, 227, 229, 229, 231, 230, 231, 230, 229, 229, 228, 229, 229, 229, 232, 232, 234, 232, 232, 228, 213, 174, 97, 93, 76, 95, 97, 131, 186, 213, 226, 229, 229, 229, 229, 228, 228, 227, 226, 228, 228, 226, 228, 230, 229, 229, 228, 228, 230, 229, 228, 228, 228, 230, 229, 228, 228, 228, 228, 230, 229, 228, 228, 228, 229, 229, 229, 226, 224, 225, 228, 227, 225, 225, 224, 226, 226, 224, 225, 224, 220, 224, 226, 225, 222, 219, 213, 213, 213, 211, 212, 215, 140, 213, 214, 217, 218, 214, 212, 212, 214, 214, 213, 216, 214, 216, 218, 217, 216, 219, 222, 222, 220, 217, 217, 219, 218, 219, 220, 224, 223, 225, 223, 225, 224, 224, 226, 225, 227, 223, 226, 227, 228, 227, 227, 226, 225, 223, 227, 226, 224, 226, 226, 228, 229, 228, 228, 227, 226, 227, 229, 227, 228, 228, 227, 228, 229, 228, 227, 229, 229, 228, 227, 227, 227, 228, 227, 228, 227, 226, 227, 227, 228, 229, 227, 227, 228, 228, 230, 228, 227, 226, 229, 228, 229, 228, 228, 230, 230, 230, 229, 228, 228, 229, 230, 229, 230, 229, 230, 230, 230, 229, 229, 229, 230, 230, 230, 228, 228, 229, 229, 230, 227, 228, 229, 231, 230, 229, 229, 230, 231, 231, 231, 230, 230, 229, 231, 231, 231, 231, 230, 230, 233, 232, 231, 231, 230, 231, 232, 232, 233, 233, 233, 232, 225, 211, 141, 77, 130, 220, 217, 197, 121, 98, 168, 219, 228, 229, 227, 229, 229, 230, 228, 228, 229, 229, 228, 229, 230, 228, 230, 231, 232, 231, 232, 232, 229, 221, 181, 109, 107, 92, 122, 109, 126, 195, 222, 227, 229, 229, 228, 228, 228, 226, 228, 228, 226, 227, 228, 228, 230, 228, 228, 228, 229, 229, 230, 228, 227, 230, 230, 230, 229, 227, 228, 230, 230, 228, 228, 227, 229, 228, 228, 227, 226, 226, 229, 227, 225, 224, 225, 226, 227, 224, 224, 221, 224, 225, 224, 227, 225, 220, 213, 215, 218, 211, 212, 215, 126, 211, 216, 218, 215, 214, 215, 212, 214, 216, 213, 215, 215, 218, 217, 218, 216, 218, 221, 224, 221, 219, 217, 221, 219, 220, 220, 222, 222, 224, 224, 223, 224, 223, 224, 224, 226, 222, 225, 225, 225, 227, 227, 226, 225, 225, 228, 226, 226, 227, 229, 228, 229, 229, 227, 226, 228, 228, 228, 227, 228, 227, 228, 228, 228, 227, 228, 228, 230, 229, 230, 228, 228, 229, 228, 227, 227, 227, 228, 226, 229, 228, 227, 227, 228, 228, 229, 228, 229, 228, 228, 229, 229, 228, 228, 229, 230, 230, 229, 228, 228, 229, 230, 230, 229, 229, 229, 229, 230, 229, 229, 229, 230, 231, 230, 229, 229, 230, 231, 230, 229, 228, 230, 230, 231, 231, 229, 230, 230, 231, 231, 230, 230, 229, 231, 232, 231, 231, 231, 232, 233, 232, 232, 232, 231, 232, 232, 233, 233, 233, 233, 230, 222, 209, 93, 78, 193, 222, 213, 168, 97, 123, 203, 226, 226, 227, 227, 230, 230, 230, 228, 226, 229, 229, 230, 230, 228, 228, 229, 231, 231, 231, 231, 231, 233, 229, 219, 173, 135, 101, 143, 126, 96, 152, 212, 227, 228, 229, 229, 228, 229, 228, 229, 228, 227, 226, 229, 229, 230, 229, 229, 228, 231, 229, 230, 228, 228, 230, 230, 231, 228, 228, 230, 230, 229, 228, 228, 228, 229, 228, 227, 226, 225, 224, 227, 229, 228, 225, 226, 227, 225, 224, 225, 221, 221, 224, 225, 226, 224, 221, 213, 217, 219, 216, 215, 217, 121, 211, 217, 218, 214, 215, 216, 218, 214, 218, 216, 219, 217, 216, 219, 220, 219, 220, 224, 224, 224, 222, 221, 221, 220, 221, 219, 224, 221, 225, 223, 224, 222, 222, 224, 222, 225, 223, 224, 224, 226, 227, 227, 226, 227, 227, 227, 228, 227, 227, 228, 230, 229, 229, 227, 227, 229, 230, 228, 228, 227, 226, 227, 229, 228, 228, 227, 229, 229, 230, 230, 229, 228, 227, 228, 227, 226, 228, 227, 228, 226, 228, 227, 227, 228, 228, 228, 228, 228, 228, 229, 229, 229, 229, 229, 230, 230, 230, 228, 228, 229, 229, 229, 229, 229, 229, 229, 230, 230, 228, 229, 229, 230, 231, 230, 230, 229, 229, 231, 230, 228, 229, 229, 230, 231, 231, 230, 231, 231, 232, 232, 229, 228, 230, 230, 231, 230, 230, 231, 231, 233, 232, 232, 231, 231, 232, 233, 233, 231, 232, 232, 228, 219, 196, 94, 102, 216, 221, 211, 133, 94, 157, 218, 228, 227, 228, 228, 230, 230, 229, 226, 228, 227, 230, 229, 229, 228, 228, 229, 229, 228, 231, 232, 231, 232, 229, 227, 216, 137, 170, 114, 163, 107, 99, 189, 224, 229, 230, 228, 227, 229, 229, 229, 229, 227, 228, 229, 229, 229, 229, 229, 228, 231, 229, 229, 228, 228, 229, 230, 230, 227, 229, 229, 230, 229, 228, 229, 228, 228, 228, 227, 227, 226, 224, 226, 228, 228, 226, 227, 227, 226, 226, 224, 221, 222, 225, 225, 225, 223, 221, 218, 218, 216, 214, 214, 219, 132, 213, 219, 220, 217, 215, 217, 217, 213, 216, 216, 215, 220, 217, 220, 221, 219, 219, 224, 225, 220, 220, 221, 220, 220, 221, 219, 221, 222, 225, 223, 225, 223, 224, 225, 223, 224, 223, 225, 225, 227, 228, 226, 226, 224, 225, 226, 226, 226, 227, 228, 229, 229, 229, 228, 227, 227, 228, 229, 229, 227, 228, 227, 229, 230, 228, 227, 229, 230, 229, 227, 228, 228, 228, 229, 229, 227, 226, 228, 228, 228, 228, 227, 227, 229, 229, 229, 229, 229, 228, 230, 230, 230, 228, 228, 230, 230, 231, 230, 229, 228, 230, 229, 229, 229, 229, 229, 230, 231, 229, 229, 230, 231, 231, 230, 229, 230, 229, 229, 229, 229, 229, 229, 230, 231, 231, 230, 230, 231, 232, 232, 230, 229, 229, 230, 231, 231, 230, 231, 232, 233, 233, 232, 231, 232, 232, 232, 233, 232, 232, 231, 227, 219, 175, 119, 136, 223, 219, 199, 108, 92, 184, 224, 227, 228, 227, 227, 229, 230, 229, 228, 226, 226, 226, 229, 229, 228, 226, 229, 230, 228, 230, 228, 231, 231, 230, 230, 221, 203, 186, 159, 178, 142, 81, 140, 216, 228, 229, 228, 228, 228, 229, 230, 229, 227, 228, 230, 231, 230, 229, 229, 229, 230, 229, 226, 228, 229, 229, 230, 231, 228, 228, 228, 230, 229, 230, 229, 229, 229, 229, 226, 226, 227, 226, 228, 228, 229, 227, 227, 227, 224, 225, 224, 221, 220, 223, 225, 226, 224, 221, 217, 218, 216, 216, 213, 218, 124, 215, 220, 221, 217, 215, 214, 217, 215, 214, 215, 215, 219, 218, 219, 220, 220, 221, 223, 224, 222, 219, 218, 220, 221, 224, 222, 220, 222, 225, 224, 224, 222, 221, 224, 223, 225, 223, 226, 225, 228, 228, 227, 224, 226, 224, 228, 226, 228, 227, 228, 228, 230, 229, 228, 228, 228, 229, 229, 227, 226, 228, 229, 229, 230, 229, 228, 229, 230, 230, 229, 227, 228, 228, 229, 229, 228, 228, 228, 228, 228, 228, 227, 227, 227, 229, 229, 227, 228, 228, 230, 230, 229, 228, 228, 230, 229, 230, 229, 229, 228, 230, 230, 229, 229, 229, 229, 230, 229, 229, 229, 229, 231, 231, 230, 229, 229, 229, 230, 230, 230, 230, 229, 230, 231, 231, 230, 231, 230, 232, 231, 230, 229, 230, 231, 231, 232, 230, 231, 231, 233, 233, 232, 231, 232, 233, 232, 233, 232, 232, 230, 227, 219, 166, 116, 159, 224, 217, 190, 99, 102, 202, 226, 228, 228, 226, 225, 227, 229, 227, 227, 227, 225, 226, 229, 229, 228, 227, 229, 230, 230, 228, 230, 230, 231, 230, 230, 227, 224, 180, 220, 157, 174, 95, 101, 205, 228, 228, 229, 229, 227, 228, 230, 227, 228, 228, 229, 230, 230, 228, 228, 229, 230, 229, 228, 229, 228, 230, 230, 230, 228, 228, 229, 231, 230, 229, 228, 228, 230, 229, 228, 225, 225, 226, 227, 227, 227, 228, 227, 228, 228, 227, 224, 222, 224, 224, 227, 226, 224, 221, 215, 217, 218, 217, 213, 219, 119, 213, 219, 221, 218, 217, 213, 216, 217, 215, 216, 216, 218, 221, 220, 220, 222, 222, 224, 221, 223, 222, 218, 218, 220, 222, 223, 221, 223, 224, 224, 221, 223, 222, 224, 225, 226, 224, 224, 225, 228, 227, 228, 225, 226, 227, 227, 228, 226, 226, 228, 230, 229, 230, 229, 227, 228, 229, 228, 227, 227, 227, 229, 229, 230, 229, 228, 229, 230, 229, 229, 227, 228, 227, 230, 229, 229, 228, 228, 230, 229, 230, 228, 228, 228, 230, 230, 229, 229, 229, 229, 230, 229, 229, 228, 229, 229, 229, 229, 229, 228, 230, 230, 229, 229, 229, 228, 229, 230, 230, 229, 229, 230, 231, 230, 230, 229, 230, 231, 231, 230, 229, 229, 230, 230, 230, 230, 230, 231, 232, 231, 230, 229, 230, 231, 231, 231, 229, 231, 231, 233, 232, 231, 230, 232, 233, 233, 233, 231, 231, 230, 228, 219, 152, 119, 178, 223, 214, 175, 93, 122, 211, 228, 226, 227, 228, 227, 226, 229, 228, 227, 228, 225, 227, 230, 229, 229, 230, 229, 230, 229, 228, 230, 230, 230, 231, 228, 229, 226, 193, 226, 166, 193, 116, 79, 180, 226, 228, 225, 227, 228, 228, 229, 227, 229, 229, 230, 229, 230, 229, 228, 229, 230, 229, 229, 229, 229, 229, 229, 230, 229, 228, 230, 230, 230, 229, 227, 229, 230, 230, 229, 225, 224, 226, 228, 228, 227, 229, 228, 228, 227, 226, 225, 223, 226, 226, 227, 226, 226, 223, 216, 216, 217, 216, 212, 218, 118, 214, 218, 220, 215, 218, 216, 215, 221, 216, 215, 217, 219, 221, 221, 222, 224, 225, 220, 224, 222, 224, 218, 221, 224, 223, 223, 221, 224, 224, 224, 223, 223, 223, 224, 223, 225, 223, 223, 226, 226, 228, 228, 225, 227, 227, 227, 228, 226, 226, 228, 230, 230, 229, 228, 227, 229, 230, 228, 228, 228, 228, 229, 230, 230, 228, 228, 230, 229, 229, 229, 228, 228, 228, 229, 228, 228, 228, 228, 230, 230, 230, 228, 228, 229, 230, 228, 228, 229, 229, 229, 230, 230, 229, 228, 229, 229, 229, 229, 229, 229, 230, 230, 229, 229, 229, 230, 230, 230, 230, 230, 230, 230, 230, 230, 230, 229, 230, 230, 231, 228, 229, 229, 230, 230, 230, 229, 230, 231, 232, 231, 230, 229, 229, 231, 231, 232, 230, 231, 232, 232, 232, 231, 231, 231, 232, 233, 232, 232, 232, 230, 226, 223, 146, 129, 193, 224, 213, 163, 93, 135, 217, 228, 226, 226, 226, 226, 227, 228, 228, 227, 227, 226, 229, 230, 229, 230, 230, 230, 230, 229, 229, 229, 230, 230, 230, 229, 230, 223, 206, 214, 167, 197, 147, 78, 156, 223, 229, 226, 226, 227, 229, 229, 228, 228, 229, 230, 231, 230, 228, 228, 229, 231, 231, 230, 229, 230, 229, 230, 230, 229, 229, 229, 231, 230, 230, 230, 228, 230, 230, 229, 225, 226, 226, 228, 228, 228, 229, 227, 227, 228, 226, 225, 225, 225, 227, 225, 225, 227, 223, 215, 211, 218, 214, 214, 216, 135, 215, 217, 217, 216, 215, 215, 218, 215, 216, 216, 219, 223, 223, 223, 221, 221, 222, 221, 221, 222, 221, 223, 223, 224, 222, 223, 223, 222, 225, 224, 223, 221, 221, 224, 222, 223, 222, 224, 227, 227, 227, 228, 226, 226, 226, 228, 228, 228, 227, 228, 230, 230, 229, 228, 228, 227, 230, 230, 229, 228, 228, 230, 230, 230, 229, 229, 230, 230, 230, 229, 228, 228, 228, 227, 229, 229, 228, 228, 230, 229, 229, 229, 228, 229, 230, 229, 228, 228, 228, 229, 230, 230, 229, 229, 230, 230, 230, 229, 229, 229, 231, 230, 230, 229, 230, 229, 230, 230, 229, 229, 230, 230, 230, 230, 230, 229, 230, 230, 231, 229, 229, 229, 230, 229, 230, 230, 230, 230, 231, 232, 231, 230, 231, 231, 230, 231, 230, 231, 232, 232, 232, 231, 231, 231, 232, 232, 232, 230, 231, 230, 224, 222, 139, 126, 201, 221, 214, 152, 85, 148, 219, 228, 228, 227, 227, 225, 228, 227, 227, 229, 226, 226, 229, 229, 229, 230, 230, 229, 230, 230, 229, 229, 229, 230, 228, 230, 230, 221, 219, 179, 165, 189, 169, 75, 124, 214, 227, 225, 226, 226, 229, 226, 225, 229, 229, 230, 230, 230, 229, 228, 228, 230, 230, 230, 229, 230, 230, 231, 231, 229, 229, 229, 230, 230, 230, 229, 229, 230, 230, 228, 227, 226, 226, 228, 228, 230, 227, 228, 227, 229, 229, 227, 227, 227, 228, 226, 225, 227, 222, 216, 213, 218, 218, 212, 219, 133, 215, 216, 215, 214, 213, 213, 215, 220, 217, 216, 220, 223, 223, 224, 223, 221, 221, 223, 222, 222, 222, 222, 222, 219, 224, 221, 223, 223, 226, 222, 223, 222, 220, 224, 220, 222, 223, 224, 227, 228, 227, 229, 228, 228, 225, 227, 228, 228, 227, 228, 229, 231, 229, 228, 228, 228, 230, 229, 228, 229, 227, 230, 229, 229, 228, 229, 230, 230, 230, 229, 228, 228, 228, 230, 229, 228, 227, 229, 229, 230, 229, 228, 228, 229, 229, 229, 228, 229, 229, 230, 231, 230, 229, 228, 230, 229, 229, 229, 229, 229, 231, 231, 230, 229, 229, 229, 230, 230, 229, 228, 229, 230, 230, 230, 229, 229, 229, 231, 231, 229, 229, 230, 230, 230, 230, 230, 230, 230, 230, 230, 230, 230, 230, 231, 231, 231, 230, 230, 232, 232, 233, 232, 231, 231, 231, 232, 232, 231, 230, 229, 224, 221, 135, 119, 202, 222, 214, 145, 85, 152, 219, 228, 230, 226, 227, 227, 228, 227, 229, 229, 229, 227, 229, 230, 231, 229, 228, 229, 230, 230, 230, 229, 228, 227, 229, 229, 228, 223, 226, 169, 191, 180, 185, 84, 104, 212, 228, 225, 225, 227, 229, 225, 227, 228, 229, 231, 230, 230, 229, 227, 230, 230, 231, 230, 230, 230, 230, 229, 231, 228, 228, 229, 230, 229, 229, 227, 229, 229, 229, 229, 228, 229, 227, 229, 227, 229, 228, 229, 228, 230, 229, 228, 227, 226, 226, 228, 226, 228, 223, 214, 214, 218, 215, 212, 220, 136, 215, 218, 216, 215, 214, 216, 216, 220, 219, 218, 218, 223, 222, 224, 222, 221, 223, 222, 222, 223, 224, 222, 223, 220, 224, 225, 223, 223, 226, 224, 224, 224, 221, 224, 221, 222, 223, 224, 227, 226, 228, 229, 227, 227, 226, 228, 230, 229, 228, 229, 229, 230, 229, 229, 228, 228, 228, 229, 229, 228, 229, 230, 229, 229, 229, 229, 229, 230, 230, 229, 229, 228, 229, 230, 229, 228, 227, 229, 230, 229, 229, 228, 228, 229, 230, 230, 229, 229, 229, 230, 231, 230, 229, 229, 229, 230, 230, 229, 229, 229, 230, 230, 230, 230, 230, 230, 230, 230, 229, 229, 228, 231, 230, 230, 229, 230, 230, 230, 231, 229, 229, 229, 230, 231, 230, 229, 230, 230, 230, 231, 231, 230, 230, 232, 232, 231, 231, 231, 232, 232, 233, 232, 232, 230, 229, 223, 228, 231, 231, 228, 223, 212, 122, 108, 213, 219, 210, 142, 81, 166, 222, 228, 229, 226, 228, 227, 228, 228, 228, 228, 228, 225, 229, 230, 230, 230, 230, 230, 230, 231, 229, 229, 227, 228, 225, 229, 226, 227, 226, 166, 202, 168, 191, 97, 94, 205, 226, 225, 224, 224, 226, 228, 227, 227, 227, 229, 231, 231, 229, 228, 229, 230, 230, 229, 229, 229, 230, 230, 229, 229, 229, 228, 229, 228, 230, 229, 228, 229, 229, 230, 228, 228, 229, 229, 228, 229, 227, 228, 229, 230, 228, 227, 227, 226, 227, 226, 228, 225, 223, 217, 216, 219, 215, 211, 219, 126, 215, 218, 217, 216, 215, 216, 218, 220, 219, 216, 221, 224, 222, 225, 219, 220, 223, 223, 220, 222, 222, 224, 222, 223, 225, 224, 222, 224, 228, 226, 224, 222, 222, 224, 223, 225, 225, 227, 227, 227, 228, 229, 227, 228, 228, 229, 230, 228, 229, 229, 230, 230, 229, 229, 228, 230, 230, 230, 229, 228, 229, 230, 230, 231, 228, 228, 228, 230, 231, 230, 229, 229, 229, 230, 228, 228, 227, 228, 230, 230, 229, 229, 229, 229, 230, 230, 229, 229, 229, 231, 230, 230, 229, 229, 230, 230, 230, 229, 229, 230, 230, 231, 230, 229, 229, 230, 230, 230, 228, 229, 229, 231, 231, 230, 230, 229, 230, 231, 231, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 232, 230, 230, 231, 232, 233, 232, 232, 233, 233, 234, 234, 232, 228, 223, 182, 124, 184, 229, 230, 226, 214, 178, 107, 110, 218, 219, 204, 145, 135, 162, 188, 198, 209, 216, 221, 219, 221, 225, 225, 227, 228, 229, 230, 229, 230, 230, 229, 230, 231, 231, 229, 228, 228, 228, 229, 227, 226, 226, 225, 163, 189, 162, 195, 105, 80, 200, 225, 222, 225, 224, 227, 228, 227, 228, 228, 229, 230, 230, 230, 228, 230, 230, 230, 230, 230, 229, 229, 229, 230, 228, 229, 227, 229, 229, 230, 228, 228, 227, 228, 229, 228, 228, 229, 230, 229, 229, 228, 228, 229, 230, 229, 228, 227, 227, 229, 227, 226, 225, 223, 218, 216, 218, 219, 215, 221, 131, 215, 220, 215, 216, 217, 217, 217, 222, 220, 219, 220, 221, 223, 224, 219, 222, 221, 222, 222, 222, 221, 226, 223, 224, 224, 221, 224, 223, 228, 227, 227, 224, 224, 225, 223, 225, 224, 225, 227, 228, 228, 228, 228, 228, 227, 230, 230, 229, 228, 229, 230, 230, 231, 229, 229, 229, 229, 230, 229, 228, 229, 230, 230, 229, 228, 229, 230, 231, 230, 229, 227, 227, 229, 229, 229, 228, 228, 229, 230, 230, 229, 228, 229, 230, 230, 230, 229, 228, 229, 230, 231, 230, 229, 229, 230, 230, 230, 229, 229, 230, 231, 231, 230, 230, 229, 230, 231, 231, 229, 229, 229, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 232, 231, 231, 231, 231, 232, 232, 231, 231, 231, 233, 234, 233, 233, 234, 235, 235, 236, 232, 228, 221, 128, 129, 113, 223, 226, 213, 175, 119, 92, 151, 203, 185, 160, 148, 147, 136, 140, 136, 137, 146, 170, 179, 183, 193, 199, 210, 222, 227, 228, 229, 229, 230, 230, 229, 231, 231, 229, 226, 223, 219, 214, 213, 213, 217, 216, 173, 208, 146, 194, 110, 76, 183, 222, 225, 226, 227, 227, 228, 226, 228, 229, 230, 229, 229, 228, 228, 229, 230, 231, 230, 230, 230, 230, 230, 230, 229, 230, 223, 229, 230, 229, 228, 229, 228, 229, 229, 228, 227, 228, 229, 229, 229, 228, 228, 228, 230, 228, 228, 228, 227, 227, 227, 226, 227, 223, 221, 220, 216, 215, 214, 220, 133, 214, 219, 216, 221, 213, 219, 218, 219, 222, 221, 220, 221, 220, 223, 223, 222, 221, 221, 221, 221, 224, 225, 221, 223, 226, 223, 225, 225, 226, 226, 226, 224, 224, 225, 224, 226, 226, 225, 227, 229, 229, 227, 227, 227, 227, 230, 229, 229, 226, 229, 230, 230, 231, 229, 229, 230, 229, 230, 229, 228, 228, 230, 230, 230, 229, 229, 229, 230, 230, 229, 229, 228, 229, 229, 229, 229, 229, 228, 230, 230, 229, 228, 229, 230, 230, 230, 229, 229, 229, 230, 231, 230, 229, 230, 230, 230, 230, 229, 229, 230, 231, 231, 230, 230, 229, 230, 231, 231, 230, 230, 230, 230, 231, 230, 230, 229, 230, 232, 230, 231, 231, 231, 232, 232, 232, 232, 231, 231, 232, 232, 231, 232, 232, 233, 234, 234, 234, 234, 235, 237, 237, 235, 231, 222, 172, 111, 113, 193, 215, 197, 139, 100, 103, 132, 139, 130, 133, 130, 134, 120, 120, 124, 115, 115, 118, 132, 137, 116, 131, 154, 189, 212, 224, 231, 230, 232, 232, 233, 232, 230, 217, 191, 173, 155, 150, 143, 135, 140, 139, 126, 198, 121, 164, 91, 104, 168, 219, 223, 224, 227, 227, 227, 227, 228, 227, 229, 229, 229, 228, 227, 228, 230, 231, 229, 229, 230, 231, 231, 231, 230, 229, 227, 230, 231, 229, 229, 229, 229, 230, 230, 229, 228, 229, 230, 229, 230, 229, 228, 229, 229, 226, 228, 227, 228, 229, 226, 226, 225, 221, 220, 220, 217, 215, 212, 218, 124, 214, 219, 220, 216, 219, 219, 223, 218, 222, 220, 220, 221, 224, 224, 221, 223, 223, 224, 221, 221, 223, 224, 218, 224, 226, 223, 224, 225, 227, 227, 226, 224, 225, 224, 225, 226, 225, 226, 227, 228, 229, 228, 228, 228, 229, 230, 230, 227, 227, 229, 230, 230, 228, 230, 228, 229, 229, 230, 229, 229, 229, 230, 231, 230, 229, 229, 230, 231, 230, 229, 229, 228, 229, 230, 230, 228, 228, 229, 230, 230, 229, 229, 229, 230, 230, 229, 229, 230, 230, 230, 231, 230, 230, 229, 230, 230, 230, 229, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 229, 231, 231, 231, 231, 230, 231, 232, 232, 232, 231, 231, 231, 232, 233, 233, 232, 232, 234, 235, 234, 234, 234, 235, 237, 237, 237, 235, 231, 222, 148, 135, 107, 137, 127, 99, 125, 134, 131, 127, 126, 124, 123, 128, 127, 124, 129, 130, 123, 122, 116, 128, 120, 83, 87, 113, 163, 199, 227, 232, 232, 232, 231, 224, 197, 168, 155, 153, 141, 145, 139, 134, 137, 134, 129, 127, 117, 120, 111, 101, 114, 173, 158, 186, 220, 216, 214, 225, 229, 228, 229, 229, 229, 228, 227, 229, 229, 230, 229, 228, 230, 230, 230, 231, 229, 229, 230, 231, 231, 230, 230, 230, 230, 230, 230, 229, 229, 228, 230, 230, 228, 228, 228, 228, 229, 228, 227, 226, 227, 226, 226, 225, 224, 220, 219, 218, 220, 216, 216, 217, 122, 210, 217, 221, 220, 217, 217, 219, 216, 220, 222, 219, 224, 222, 224, 222, 221, 224, 222, 222, 224, 223, 224, 222, 221, 224, 223, 222, 225, 228, 227, 226, 226, 225, 226, 227, 228, 225, 225, 226, 228, 228, 229, 229, 229, 228, 231, 230, 227, 228, 230, 231, 231, 230, 230, 229, 228, 229, 231, 230, 229, 230, 230, 230, 230, 230, 229, 229, 230, 230, 229, 229, 229, 229, 229, 230, 228, 229, 229, 229, 229, 229, 229, 229, 230, 230, 229, 229, 229, 229, 230, 230, 230, 229, 229, 230, 230, 231, 230, 230, 229, 231, 231, 230, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 231, 231, 230, 232, 232, 232, 231, 231, 231, 232, 232, 232, 232, 232, 233, 234, 234, 234, 234, 234, 235, 237, 237, 234, 232, 227, 159, 156, 123, 99, 123, 133, 139, 145, 140, 138, 142, 136, 142, 136, 138, 140, 142, 134, 131, 122, 122, 124, 128, 103, 64, 67, 93, 147, 202, 229, 231, 228, 221, 185, 162, 162, 156, 162, 161, 160, 162, 152, 155, 147, 149, 137, 127, 117, 114, 125, 128, 107, 128, 86, 163, 132, 131, 199, 226, 228, 228, 229, 229, 228, 227, 230, 230, 230, 229, 230, 230, 230, 231, 230, 229, 230, 229, 230, 231, 231, 230, 229, 230, 231, 230, 228, 228, 228, 230, 230, 228, 227, 228, 226, 228, 226, 227, 225, 223, 226, 225, 223, 223, 220, 217, 218, 220, 219, 212, 218, 116, 211, 217, 218, 218, 217, 217, 216, 218, 217, 220, 218, 221, 224, 223, 222, 220, 223, 220, 224, 226, 224, 223, 222, 221, 223, 222, 223, 223, 226, 227, 226, 225, 226, 224, 227, 225, 226, 227, 227, 227, 228, 229, 228, 229, 230, 231, 230, 228, 229, 230, 230, 231, 230, 230, 229, 230, 229, 230, 229, 229, 228, 230, 230, 230, 229, 229, 230, 230, 230, 230, 229, 228, 228, 229, 227, 229, 229, 229, 229, 229, 229, 228, 229, 230, 230, 230, 229, 229, 228, 229, 230, 230, 229, 229, 230, 230, 230, 230, 230, 229, 230, 231, 231, 229, 230, 230, 231, 231, 230, 230, 229, 231, 231, 231, 230, 231, 231, 232, 232, 231, 231, 231, 231, 233, 231, 230, 231, 231, 232, 233, 233, 232, 232, 233, 234, 234, 234, 234, 235, 235, 236, 236, 234, 230, 222, 163, 130, 111, 133, 135, 141, 148, 145, 139, 137, 144, 143, 148, 148, 145, 148, 147, 146, 141, 133, 131, 127, 124, 130, 77, 70, 92, 104, 160, 212, 223, 219, 180, 151, 136, 135, 127, 137, 158, 160, 163, 168, 168, 164, 165, 157, 152, 142, 131, 132, 126, 128, 116, 84, 70, 64, 78, 174, 225, 227, 229, 228, 230, 227, 227, 228, 229, 230, 230, 230, 230, 231, 230, 230, 230, 229, 229, 231, 230, 231, 229, 230, 231, 230, 229, 229, 229, 229, 230, 229, 229, 227, 226, 226, 228, 229, 227, 227, 225, 228, 227, 223, 224, 218, 218, 219, 216, 218, 216, 219, 135, 213, 221, 220, 220, 218, 220, 217, 220, 218, 215, 219, 219, 224, 224, 221, 222, 223, 224, 224, 227, 226, 224, 224, 224, 226, 224, 224, 224, 227, 227, 226, 226, 225, 224, 225, 227, 226, 226, 227, 229, 229, 230, 228, 228, 229, 231, 230, 230, 228, 229, 229, 230, 231, 229, 229, 229, 230, 230, 230, 229, 228, 230, 230, 230, 229, 229, 230, 231, 230, 230, 228, 229, 229, 227, 229, 229, 228, 229, 230, 230, 230, 229, 228, 230, 230, 230, 229, 229, 228, 230, 230, 230, 229, 229, 230, 231, 231, 230, 230, 229, 231, 231, 231, 230, 229, 230, 232, 232, 231, 230, 230, 231, 231, 231, 230, 230, 231, 231, 232, 231, 231, 231, 232, 231, 232, 231, 232, 232, 233, 234, 233, 232, 232, 233, 235, 235, 235, 234, 235, 236, 237, 236, 233, 228, 213, 143, 141, 120, 119, 129, 145, 145, 147, 148, 150, 153, 153, 164, 161, 162, 160, 163, 155, 150, 144, 137, 125, 134, 129, 96, 66, 109, 86, 113, 140, 163, 157, 102, 60, 54, 54, 58, 71, 90, 106, 143, 162, 167, 174, 173, 169, 165, 158, 148, 144, 137, 128, 112, 104, 84, 57, 79, 153, 206, 221, 227, 229, 230, 228, 227, 228, 229, 230, 231, 230, 229, 230, 230, 231, 230, 229, 229, 230, 230, 231, 229, 230, 230, 229, 229, 229, 229, 229, 230, 229, 230, 229, 228, 226, 228, 226, 228, 227, 226, 226, 226, 226, 224, 219, 219, 218, 220, 219, 218, 221, 148, 215, 220, 219, 219, 219, 219, 220, 220, 221, 217, 217, 220, 222, 222, 224, 222, 223, 224, 226, 226, 227, 224, 222, 225, 226, 224, 225, 226, 224, 226, 227, 227, 225, 225, 227, 225, 228, 227, 226, 227, 229, 229, 228, 227, 228, 230, 231, 230, 228, 228, 230, 230, 230, 230, 230, 229, 231, 231, 230, 229, 230, 231, 231, 230, 229, 229, 230, 230, 231, 230, 229, 229, 229, 230, 228, 229, 228, 228, 230, 231, 230, 229, 229, 229, 231, 231, 229, 228, 229, 230, 230, 231, 229, 229, 229, 230, 230, 230, 229, 229, 231, 231, 231, 230, 229, 230, 231, 232, 231, 230, 230, 231, 231, 231, 231, 230, 231, 231, 232, 231, 230, 230, 232, 231, 231, 231, 231, 231, 232, 233, 232, 232, 232, 233, 234, 234, 234, 234, 235, 236, 236, 234, 229, 217, 190, 144, 135, 124, 130, 136, 144, 147, 154, 158, 163, 165, 169, 170, 168, 171, 169, 172, 166, 167, 158, 143, 133, 129, 86, 103, 55, 126, 92, 148, 107, 100, 85, 42, 51, 57, 63, 64, 60, 53, 53, 63, 77, 110, 155, 175, 170, 172, 177, 170, 165, 154, 150, 132, 123, 110, 111, 75, 85, 143, 188, 217, 228, 228, 227, 227, 228, 229, 231, 230, 230, 230, 230, 230, 230, 230, 229, 228, 229, 229, 230, 230, 229, 230, 230, 229, 229, 230, 229, 229, 230, 229, 227, 227, 227, 227, 227, 227, 227, 226, 228, 229, 228, 225, 224, 219, 215, 220, 219, 217, 223, 130, 215, 222, 220, 220, 221, 220, 221, 222, 221, 220, 221, 222, 224, 226, 225, 222, 223, 224, 224, 224, 225, 224, 222, 225, 225, 225, 225, 225, 225, 226, 226, 227, 226, 226, 228, 227, 227, 228, 226, 227, 229, 229, 227, 226, 228, 230, 231, 229, 229, 228, 230, 230, 230, 229, 230, 230, 231, 231, 230, 229, 230, 231, 231, 230, 229, 229, 229, 231, 231, 229, 229, 229, 230, 229, 230, 228, 228, 228, 230, 231, 230, 228, 228, 230, 230, 230, 230, 229, 229, 230, 231, 229, 229, 229, 230, 231, 231, 229, 229, 229, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 232, 231, 230, 230, 231, 232, 232, 231, 231, 232, 233, 233, 232, 232, 233, 234, 234, 234, 234, 234, 235, 236, 234, 228, 206, 174, 166, 153, 151, 143, 142, 151, 155, 152, 163, 168, 174, 173, 179, 178, 179, 176, 181, 174, 176, 172, 164, 149, 128, 90, 63, 72, 66, 67, 76, 140, 88, 159, 123, 43, 54, 76, 86, 77, 59, 58, 66, 57, 56, 78, 152, 113, 154, 174, 181, 186, 181, 173, 166, 158, 142, 123, 117, 115, 82, 66, 112, 173, 214, 223, 226, 227, 228, 229, 230, 230, 230, 230, 230, 231, 229, 229, 230, 229, 230, 230, 230, 230, 229, 229, 230, 229, 230, 230, 230, 230, 229, 229, 228, 228, 228, 229, 227, 228, 226, 227, 227, 226, 228, 228, 225, 220, 216, 221, 221, 215, 219, 137, 218, 223, 224, 221, 221, 219, 224, 221, 219, 222, 220, 223, 226, 227, 225, 225, 226, 226, 224, 223, 223, 224, 224, 227, 225, 225, 225, 224, 227, 225, 226, 227, 224, 227, 227, 228, 228, 227, 226, 228, 230, 228, 228, 227, 229, 229, 230, 229, 230, 229, 229, 230, 230, 229, 230, 230, 230, 230, 230, 229, 229, 231, 230, 230, 229, 229, 230, 231, 230, 229, 228, 229, 228, 230, 230, 229, 228, 229, 230, 230, 230, 229, 229, 230, 231, 230, 229, 229, 229, 230, 230, 230, 229, 229, 230, 231, 230, 229, 229, 230, 230, 231, 231, 230, 229, 231, 232, 231, 230, 230, 230, 232, 231, 231, 231, 230, 231, 232, 232, 231, 231, 230, 232, 232, 232, 231, 231, 232, 232, 233, 233, 232, 233, 234, 234, 235, 234, 235, 234, 233, 225, 195, 171, 157, 152, 144, 146, 146, 152, 158, 164, 169, 176, 173, 179, 184, 187, 187, 182, 182, 183, 190, 184, 180, 161, 136, 79, 54, 55, 59, 54, 64, 66, 108, 127, 87, 55, 44, 51, 76, 107, 136, 156, 149, 168, 160, 113, 162, 85, 57, 64, 112, 157, 185, 184, 181, 175, 171, 155, 148, 132, 112, 121, 75, 57, 97, 156, 208, 225, 227, 228, 230, 231, 231, 230, 230, 230, 230, 230, 225, 229, 230, 228, 231, 231, 230, 229, 229, 229, 230, 229, 229, 230, 230, 230, 230, 228, 229, 229, 229, 228, 226, 228, 227, 228, 227, 229, 226, 224, 222, 218, 222, 219, 219, 219, 150, 218, 222, 226, 220, 221, 220, 226, 223, 221, 223, 221, 223, 225, 223, 225, 226, 226, 225, 224, 225, 224, 224, 224, 224, 226, 224, 225, 226, 226, 226, 227, 225, 225, 227, 228, 229, 227, 226, 228, 230, 228, 229, 227, 226, 228, 229, 229, 228, 229, 229, 230, 231, 230, 230, 230, 230, 231, 230, 230, 230, 229, 229, 230, 230, 230, 229, 230, 231, 230, 230, 229, 229, 229, 230, 229, 228, 229, 229, 231, 230, 230, 229, 229, 230, 230, 230, 229, 230, 230, 231, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 232, 230, 230, 230, 231, 231, 232, 231, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 232, 233, 232, 233, 233, 233, 234, 235, 235, 234, 234, 230, 224, 188, 169, 156, 150, 151, 148, 155, 154, 163, 170, 178, 184, 183, 185, 187, 190, 192, 192, 188, 187, 188, 188, 184, 171, 135, 74, 57, 55, 57, 54, 63, 87, 109, 182, 210, 190, 65, 62, 71, 172, 185, 126, 144, 134, 160, 157, 139, 123, 50, 52, 53, 55, 71, 128, 171, 176, 180, 176, 166, 157, 143, 128, 123, 130, 70, 63, 93, 155, 208, 224, 229, 230, 231, 231, 230, 230, 230, 230, 229, 228, 225, 229, 226, 230, 230, 229, 229, 230, 229, 230, 229, 229, 230, 230, 230, 230, 226, 229, 229, 228, 229, 225, 228, 228, 229, 228, 228, 227, 225, 223, 221, 218, 219, 215, 222, 135, 219, 221, 224, 220, 221, 221, 222, 222, 220, 221, 221, 224, 225, 225, 225, 225, 226, 225, 224, 225, 225, 226, 225, 227, 226, 223, 225, 226, 226, 226, 227, 226, 224, 227, 229, 229, 228, 228, 228, 229, 227, 229, 228, 227, 227, 230, 230, 228, 228, 230, 231, 231, 230, 229, 229, 230, 231, 230, 229, 229, 229, 230, 230, 230, 230, 229, 230, 231, 231, 230, 229, 228, 230, 231, 228, 227, 229, 230, 231, 231, 230, 230, 230, 231, 230, 230, 229, 230, 229, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 231, 232, 231, 230, 230, 231, 232, 231, 231, 230, 231, 231, 231, 231, 230, 231, 231, 231, 231, 231, 231, 231, 232, 233, 232, 231, 231, 233, 233, 232, 233, 233, 233, 235, 234, 235, 233, 231, 223, 190, 168, 157, 150, 152, 152, 154, 162, 165, 174, 180, 188, 187, 193, 195, 195, 196, 192, 199, 196, 196, 192, 184, 171, 125, 64, 58, 58, 55, 57, 69, 97, 139, 139, 165, 182, 186, 114, 112, 146, 200, 106, 80, 60, 59, 65, 63, 61, 72, 67, 75, 66, 49, 61, 71, 86, 132, 166, 177, 179, 166, 161, 151, 130, 119, 117, 60, 70, 88, 156, 210, 226, 227, 230, 230, 229, 229, 230, 231, 230, 230, 224, 223, 230, 230, 230, 229, 229, 230, 230, 231, 229, 230, 229, 229, 229, 231, 229, 228, 230, 229, 228, 228, 229, 228, 228, 228, 228, 228, 226, 221, 219, 222, 220, 217, 222, 127, 216, 222, 223, 222, 222, 223, 222, 222, 219, 222, 219, 223, 225, 225, 224, 224, 225, 227, 225, 225, 224, 225, 224, 224, 226, 226, 227, 226, 226, 227, 227, 225, 225, 228, 228, 229, 228, 228, 229, 230, 230, 229, 228, 228, 229, 229, 230, 229, 229, 229, 231, 231, 230, 230, 229, 230, 231, 231, 229, 228, 229, 230, 230, 231, 230, 229, 230, 230, 230, 230, 228, 228, 230, 230, 229, 229, 229, 229, 230, 230, 230, 229, 229, 231, 230, 231, 229, 229, 230, 231, 231, 230, 230, 230, 230, 230, 231, 229, 229, 230, 231, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 231, 231, 230, 231, 231, 231, 231, 231, 232, 233, 232, 232, 232, 232, 232, 233, 233, 232, 233, 232, 235, 234, 234, 230, 225, 193, 168, 163, 156, 150, 152, 157, 165, 166, 174, 179, 185, 192, 195, 204, 200, 202, 201, 197, 201, 196, 191, 182, 156, 101, 68, 105, 153, 128, 99, 95, 107, 135, 134, 136, 143, 135, 142, 137, 136, 140, 139, 133, 125, 114, 105, 89, 71, 67, 69, 69, 79, 73, 67, 61, 55, 59, 56, 85, 151, 176, 173, 171, 163, 142, 123, 127, 110, 56, 60, 97, 175, 220, 228, 230, 229, 229, 229, 230, 232, 229, 229, 229, 230, 231, 230, 230, 229, 230, 231, 231, 231, 230, 229, 229, 231, 230, 230, 229, 228, 230, 231, 228, 228, 228, 225, 228, 230, 228, 227, 225, 221, 219, 222, 217, 217, 222, 126, 216, 222, 221, 220, 221, 221, 221, 221, 220, 220, 220, 222, 224, 225, 225, 222, 225, 226, 226, 227, 225, 226, 226, 224, 226, 226, 226, 226, 227, 228, 228, 225, 227, 228, 229, 230, 228, 227, 228, 229, 230, 230, 228, 227, 228, 229, 230, 229, 229, 230, 230, 230, 230, 229, 229, 230, 230, 230, 230, 228, 229, 230, 230, 231, 230, 230, 230, 231, 230, 229, 229, 229, 231, 231, 230, 229, 229, 229, 230, 230, 230, 230, 230, 230, 230, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 229, 229, 230, 231, 232, 231, 230, 229, 230, 231, 232, 230, 230, 230, 231, 231, 232, 230, 231, 231, 232, 232, 232, 231, 230, 232, 233, 233, 232, 231, 232, 233, 234, 232, 232, 234, 235, 234, 233, 228, 204, 169, 165, 160, 162, 159, 159, 164, 172, 176, 180, 185, 188, 200, 203, 208, 202, 207, 201, 203, 204, 193, 180, 145, 73, 60, 62, 86, 107, 100, 117, 131, 140, 145, 143, 147, 147, 149, 144, 141, 147, 147, 148, 145, 144, 151, 143, 132, 121, 108, 91, 81, 81, 76, 68, 66, 55, 51, 37, 51, 70, 137, 166, 176, 164, 148, 134, 121, 133, 83, 48, 75, 118, 195, 224, 229, 230, 230, 230, 230, 231, 231, 229, 229, 229, 231, 231, 230, 230, 229, 230, 231, 231, 230, 229, 229, 230, 230, 230, 229, 229, 230, 230, 230, 228, 228, 225, 228, 228, 227, 229, 225, 222, 220, 222, 218, 218, 222, 124, 217, 223, 223, 223, 219, 220, 220, 220, 217, 222, 221, 223, 226, 225, 224, 225, 225, 226, 228, 226, 224, 225, 225, 225, 225, 225, 225, 226, 227, 229, 227, 226, 227, 226, 229, 228, 228, 228, 228, 230, 230, 229, 229, 229, 229, 230, 231, 230, 230, 229, 230, 230, 230, 230, 229, 230, 231, 230, 229, 228, 229, 231, 231, 230, 230, 230, 230, 230, 230, 230, 230, 229, 230, 231, 231, 229, 229, 230, 231, 231, 231, 229, 230, 231, 231, 230, 229, 229, 230, 231, 231, 230, 229, 230, 231, 231, 230, 229, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 232, 232, 231, 230, 231, 231, 232, 232, 231, 232, 231, 232, 233, 233, 232, 232, 232, 233, 233, 233, 233, 233, 234, 234, 231, 220, 181, 163, 158, 163, 160, 166, 165, 174, 179, 183, 191, 195, 200, 210, 208, 221, 215, 214, 205, 203, 195, 169, 106, 64, 62, 66, 88, 106, 115, 133, 148, 153, 149, 145, 144, 150, 152, 156, 162, 165, 164, 168, 167, 176, 174, 179, 180, 173, 169, 159, 146, 123, 106, 87, 60, 61, 50, 48, 43, 49, 54, 68, 117, 162, 165, 161, 148, 126, 124, 130, 55, 52, 84, 146, 211, 228, 230, 228, 229, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 229, 229, 229, 230, 230, 229, 229, 230, 230, 231, 231, 230, 228, 228, 226, 226, 229, 227, 229, 225, 222, 219, 218, 218, 217, 224, 132, 216, 221, 225, 221, 221, 218, 219, 221, 220, 222, 221, 222, 225, 226, 224, 223, 225, 225, 225, 224, 222, 223, 224, 225, 224, 225, 225, 225, 228, 227, 228, 227, 226, 226, 229, 229, 228, 227, 229, 230, 230, 230, 230, 229, 229, 229, 230, 229, 229, 230, 230, 230, 230, 229, 230, 230, 231, 230, 230, 229, 230, 231, 230, 230, 230, 230, 229, 229, 230, 230, 229, 229, 230, 231, 231, 229, 229, 230, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 230, 230, 230, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 232, 231, 231, 231, 232, 233, 233, 232, 231, 232, 233, 233, 233, 233, 232, 234, 233, 229, 195, 172, 167, 164, 167, 166, 171, 176, 181, 189, 193, 193, 202, 206, 212, 233, 234, 220, 210, 204, 184, 143, 81, 67, 70, 83, 109, 120, 128, 147, 153, 150, 148, 145, 145, 155, 163, 162, 163, 171, 186, 191, 198, 200, 208, 210, 214, 218, 219, 210, 204, 192, 178, 168, 142, 111, 71, 51, 47, 51, 55, 54, 57, 68, 91, 152, 161, 156, 136, 123, 133, 83, 51, 65, 102, 192, 227, 229, 228, 229, 229, 231, 230, 230, 229, 229, 231, 231, 230, 230, 230, 230, 231, 230, 229, 228, 228, 231, 230, 230, 229, 230, 231, 231, 231, 229, 227, 226, 225, 228, 227, 229, 225, 224, 219, 220, 218, 218, 221, 138, 219, 224, 224, 221, 223, 220, 220, 220, 221, 222, 221, 225, 223, 224, 224, 224, 224, 225, 226, 223, 224, 224, 224, 225, 225, 226, 224, 226, 227, 226, 228, 227, 226, 227, 228, 228, 227, 228, 228, 229, 229, 229, 230, 228, 229, 230, 230, 229, 229, 230, 230, 230, 230, 229, 230, 229, 230, 230, 229, 229, 229, 230, 231, 230, 229, 229, 230, 230, 230, 230, 229, 229, 230, 230, 230, 229, 230, 230, 231, 230, 229, 229, 229, 230, 231, 231, 230, 230, 230, 230, 230, 230, 229, 230, 230, 231, 231, 229, 229, 229, 230, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 232, 232, 232, 231, 231, 230, 232, 232, 231, 231, 231, 233, 233, 233, 231, 231, 231, 234, 233, 233, 233, 233, 234, 231, 223, 182, 167, 164, 168, 168, 169, 176, 183, 188, 191, 197, 198, 205, 212, 224, 236, 234, 213, 198, 166, 105, 61, 60, 75, 108, 122, 133, 142, 150, 156, 148, 140, 147, 155, 160, 161, 166, 180, 189, 195, 200, 201, 204, 207, 206, 210, 217, 220, 226, 227, 229, 229, 225, 214, 195, 173, 150, 111, 67, 53, 57, 59, 61, 68, 65, 87, 145, 150, 149, 131, 124, 124, 48, 60, 74, 165, 220, 229, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 229, 230, 231, 231, 229, 227, 228, 229, 230, 230, 229, 230, 230, 230, 230, 229, 227, 226, 224, 226, 230, 228, 225, 223, 219, 220, 218, 216, 219, 124, 217, 224, 221, 223, 222, 222, 223, 224, 221, 222, 220, 223, 226, 224, 225, 226, 224, 225, 228, 225, 224, 224, 225, 225, 224, 224, 225, 225, 229, 226, 228, 227, 226, 228, 228, 228, 228, 228, 227, 229, 229, 230, 229, 228, 229, 230, 231, 229, 229, 229, 230, 231, 231, 230, 229, 228, 230, 229, 229, 228, 230, 231, 230, 230, 229, 230, 230, 230, 230, 230, 229, 229, 230, 231, 231, 229, 230, 229, 230, 230, 231, 230, 230, 230, 231, 231, 229, 230, 230, 231, 231, 230, 229, 229, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 230, 230, 230, 231, 232, 232, 231, 231, 231, 232, 233, 231, 231, 231, 233, 233, 232, 231, 231, 232, 233, 233, 233, 233, 232, 233, 229, 213, 175, 166, 167, 170, 173, 177, 181, 189, 186, 193, 199, 202, 210, 216, 221, 232, 220, 189, 125, 60, 53, 66, 99, 117, 126, 137, 152, 159, 154, 142, 142, 159, 160, 152, 156, 169, 178, 185, 194, 200, 196, 199, 202, 205, 207, 209, 213, 220, 224, 223, 226, 226, 229, 233, 232, 223, 205, 171, 145, 104, 54, 50, 62, 64, 68, 70, 84, 145, 144, 141, 121, 143, 55, 52, 81, 133, 214, 229, 228, 230, 231, 231, 232, 230, 230, 230, 231, 229, 231, 230, 229, 230, 230, 231, 230, 227, 227, 229, 230, 231, 229, 230, 230, 231, 229, 230, 228, 229, 226, 227, 230, 227, 222, 222, 218, 221, 222, 218, 217, 143, 217, 223, 224, 224, 222, 222, 223, 222, 223, 221, 221, 223, 225, 226, 225, 225, 226, 224, 227, 226, 222, 224, 224, 225, 224, 222, 224, 224, 226, 226, 229, 227, 227, 227, 229, 229, 229, 228, 228, 229, 230, 230, 228, 228, 230, 230, 230, 229, 229, 230, 231, 231, 231, 229, 229, 229, 229, 229, 229, 229, 230, 231, 230, 231, 229, 230, 230, 230, 230, 230, 229, 229, 230, 231, 230, 229, 229, 230, 230, 230, 230, 230, 230, 230, 231, 231, 229, 230, 230, 231, 231, 230, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 232, 230, 230, 230, 231, 232, 232, 231, 230, 232, 232, 232, 231, 231, 231, 232, 232, 233, 231, 232, 232, 234, 234, 234, 233, 233, 232, 229, 203, 174, 171, 172, 176, 177, 178, 186, 187, 193, 195, 203, 211, 209, 217, 213, 208, 166, 79, 64, 67, 88, 104, 121, 126, 147, 158, 156, 150, 142, 150, 165, 156, 152, 155, 174, 177, 178, 169, 161, 151, 141, 140, 143, 148, 157, 171, 187, 206, 219, 223, 223, 226, 228, 228, 233, 232, 233, 224, 201, 168, 132, 77, 56, 55, 61, 68, 71, 99, 141, 142, 135, 137, 70, 52, 70, 108, 204, 228, 229, 228, 230, 232, 231, 230, 230, 230, 231, 231, 230, 229, 229, 230, 231, 230, 230, 228, 228, 229, 230, 229, 229, 230, 230, 231, 229, 228, 228, 228, 226, 227, 227, 226, 224, 223, 218, 221, 221, 216, 219, 123, 214, 225, 224, 223, 220, 220, 226, 226, 222, 220, 222, 224, 225, 226, 226, 225, 224, 227, 227, 225, 224, 223, 227, 225, 225, 223, 224, 223, 227, 227, 227, 226, 228, 228, 228, 229, 228, 228, 228, 229, 230, 230, 229, 229, 230, 230, 229, 228, 228, 229, 230, 230, 231, 229, 228, 229, 230, 229, 229, 229, 229, 230, 231, 231, 230, 230, 230, 230, 230, 230, 230, 229, 230, 231, 230, 229, 229, 230, 231, 230, 230, 230, 230, 230, 231, 231, 229, 230, 230, 231, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 231, 232, 232, 232, 231, 231, 232, 232, 232, 232, 232, 231, 232, 233, 233, 231, 232, 233, 233, 234, 234, 233, 233, 233, 230, 202, 180, 178, 180, 179, 185, 184, 193, 193, 201, 205, 207, 212, 208, 197, 170, 118, 66, 69, 104, 95, 106, 122, 129, 148, 160, 167, 158, 138, 159, 165, 155, 152, 163, 154, 144, 134, 93, 65, 54, 48, 53, 59, 106, 149, 52, 53, 68, 95, 136, 173, 201, 219, 225, 230, 228, 231, 233, 235, 234, 222, 194, 154, 106, 55, 45, 57, 62, 62, 102, 136, 144, 142, 91, 49, 65, 90, 193, 226, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 230, 230, 230, 230, 229, 229, 230, 229, 230, 229, 230, 229, 230, 230, 229, 228, 228, 228, 227, 227, 227, 225, 223, 221, 222, 216, 218, 218, 110, 212, 224, 225, 223, 222, 222, 226, 225, 224, 225, 224, 225, 226, 223, 226, 224, 224, 229, 226, 226, 223, 224, 226, 227, 228, 226, 227, 225, 226, 228, 228, 226, 227, 228, 228, 229, 228, 227, 227, 230, 230, 230, 229, 229, 229, 231, 230, 229, 229, 229, 230, 231, 230, 230, 229, 230, 231, 230, 229, 229, 229, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 230, 230, 229, 230, 229, 231, 230, 230, 229, 230, 231, 231, 231, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 231, 232, 232, 232, 231, 231, 232, 233, 233, 232, 231, 231, 232, 233, 233, 232, 232, 233, 233, 234, 234, 234, 233, 233, 231, 207, 183, 180, 182, 187, 190, 196, 197, 198, 201, 207, 208, 196, 169, 118, 67, 70, 93, 83, 107, 133, 124, 135, 153, 165, 169, 160, 145, 164, 165, 143, 148, 152, 129, 116, 78, 44, 46, 48, 55, 96, 93, 75, 89, 117, 67, 64, 68, 47, 52, 60, 81, 140, 189, 215, 227, 229, 230, 235, 237, 235, 230, 210, 170, 121, 59, 46, 50, 57, 70, 122, 146, 145, 95, 53, 68, 92, 189, 226, 228, 229, 231, 231, 231, 230, 230, 230, 232, 231, 231, 230, 230, 230, 231, 230, 229, 229, 229, 230, 231, 231, 229, 230, 229, 230, 230, 229, 228, 228, 230, 228, 227, 230, 224, 224, 222, 220, 220, 218, 221, 120, 216, 226, 222, 222, 221, 224, 226, 224, 224, 225, 225, 225, 225, 225, 225, 225, 225, 228, 227, 226, 225, 226, 226, 227, 227, 226, 227, 225, 227, 229, 227, 227, 228, 229, 230, 229, 228, 227, 228, 230, 230, 230, 228, 228, 230, 231, 230, 229, 229, 229, 230, 230, 230, 230, 228, 228, 230, 231, 230, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 230, 230, 229, 230, 231, 230, 230, 230, 230, 230, 231, 229, 230, 230, 231, 231, 231, 230, 229, 229, 231, 231, 230, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 232, 231, 230, 230, 230, 232, 232, 232, 231, 231, 232, 233, 233, 231, 231, 231, 232, 233, 233, 232, 232, 233, 234, 234, 234, 234, 234, 234, 231, 215, 180, 184, 187, 193, 196, 203, 198, 207, 200, 193, 171, 118, 75, 76, 100, 123, 123, 107, 127, 131, 138, 159, 172, 176, 157, 146, 169, 160, 145, 139, 120, 86, 59, 59, 115, 45, 40, 50, 80, 160, 163, 133, 61, 128, 121, 75, 93, 119, 78, 45, 44, 56, 76, 122, 190, 223, 230, 233, 235, 235, 236, 232, 220, 181, 134, 70, 53, 59, 70, 80, 141, 152, 84, 45, 58, 88, 194, 226, 230, 229, 231, 231, 231, 230, 229, 231, 231, 231, 231, 230, 229, 230, 231, 231, 229, 229, 230, 230, 231, 230, 228, 228, 230, 231, 230, 227, 227, 229, 230, 229, 229, 229, 224, 223, 220, 221, 224, 218, 222, 124, 213, 226, 223, 220, 218, 224, 226, 223, 225, 224, 224, 224, 227, 225, 224, 224, 225, 227, 226, 226, 225, 228, 228, 227, 227, 225, 227, 226, 228, 228, 227, 227, 227, 228, 230, 229, 227, 227, 228, 230, 229, 230, 229, 229, 230, 231, 231, 229, 229, 229, 231, 230, 230, 230, 227, 229, 231, 230, 230, 230, 230, 231, 230, 231, 230, 230, 230, 230, 231, 230, 230, 230, 230, 231, 230, 230, 229, 229, 230, 231, 231, 230, 230, 231, 231, 231, 230, 229, 229, 230, 230, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 230, 231, 232, 232, 231, 231, 232, 233, 232, 232, 231, 232, 232, 233, 233, 232, 232, 233, 234, 235, 234, 234, 235, 235, 232, 226, 191, 186, 191, 198, 205, 206, 198, 189, 162, 119, 81, 91, 117, 133, 140, 144, 138, 136, 138, 140, 159, 176, 176, 162, 145, 172, 166, 133, 127, 99, 90, 55, 47, 48, 91, 107, 43, 43, 86, 152, 169, 145, 116, 158, 62, 45, 51, 124, 151, 61, 46, 46, 45, 57, 79, 144, 206, 230, 232, 235, 236, 235, 233, 223, 187, 139, 78, 51, 55, 61, 118, 150, 62, 46, 58, 97, 200, 227, 228, 229, 231, 232, 231, 229, 230, 230, 231, 231, 231, 229, 230, 230, 231, 231, 229, 228, 230, 231, 230, 230, 228, 227, 230, 230, 230, 230, 229, 230, 230, 230, 230, 230, 226, 223, 219, 225, 222, 220, 222, 119, 214, 223, 224, 222, 218, 221, 227, 223, 225, 224, 224, 225, 225, 225, 223, 227, 225, 227, 225, 224, 224, 225, 227, 226, 227, 227, 226, 226, 229, 228, 229, 227, 227, 229, 229, 229, 227, 225, 227, 230, 230, 230, 229, 230, 230, 231, 231, 228, 229, 229, 230, 231, 229, 229, 228, 229, 231, 230, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 230, 230, 229, 229, 230, 231, 230, 230, 229, 230, 231, 230, 230, 229, 230, 231, 231, 230, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 232, 231, 230, 232, 232, 232, 231, 231, 231, 233, 233, 233, 232, 232, 233, 234, 235, 235, 234, 234, 236, 235, 230, 208, 190, 196, 197, 194, 186, 149, 106, 90, 105, 129, 137, 136, 140, 144, 141, 136, 137, 142, 162, 180, 182, 171, 142, 172, 167, 130, 110, 96, 77, 175, 68, 45, 46, 54, 120, 84, 48, 87, 141, 170, 150, 144, 160, 50, 42, 53, 86, 157, 127, 36, 38, 40, 43, 52, 80, 126, 180, 224, 232, 235, 235, 235, 234, 225, 190, 144, 76, 46, 63, 98, 145, 50, 47, 61, 126, 213, 228, 229, 229, 231, 231, 230, 229, 229, 228, 230, 230, 230, 229, 230, 230, 230, 231, 228, 229, 230, 230, 230, 229, 228, 227, 229, 230, 229, 230, 230, 229, 230, 230, 228, 230, 224, 222, 217, 225, 222, 219, 222, 111, 213, 224, 224, 221, 221, 221, 224, 221, 225, 226, 223, 225, 228, 225, 225, 227, 227, 226, 226, 225, 224, 226, 227, 226, 226, 227, 226, 224, 229, 227, 228, 228, 227, 228, 229, 230, 227, 226, 227, 229, 231, 230, 229, 229, 230, 231, 230, 229, 230, 229, 230, 230, 230, 230, 229, 229, 230, 231, 230, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 229, 230, 230, 230, 230, 229, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 231, 231, 230, 232, 232, 232, 231, 231, 231, 232, 232, 231, 231, 232, 233, 233, 233, 232, 232, 233, 234, 235, 235, 235, 235, 236, 236, 234, 224, 203, 202, 179, 148, 126, 114, 126, 146, 150, 154, 149, 141, 143, 142, 144, 141, 131, 154, 183, 186, 181, 146, 169, 174, 139, 92, 59, 62, 81, 121, 116, 98, 51, 95, 108, 147, 59, 69, 126, 167, 152, 151, 154, 45, 39, 46, 73, 150, 149, 39, 36, 39, 53, 64, 101, 164, 75, 152, 219, 233, 233, 235, 235, 234, 225, 188, 135, 68, 59, 87, 108, 46, 50, 74, 176, 225, 228, 230, 229, 230, 231, 231, 229, 229, 230, 231, 231, 230, 230, 229, 231, 230, 231, 229, 229, 229, 230, 230, 229, 227, 228, 230, 230, 231, 230, 230, 228, 230, 230, 230, 229, 224, 220, 218, 227, 219, 220, 220, 117, 213, 224, 223, 224, 225, 223, 225, 223, 223, 225, 226, 226, 228, 225, 226, 226, 225, 226, 227, 227, 225, 226, 226, 227, 227, 227, 226, 225, 228, 228, 228, 228, 226, 227, 228, 227, 227, 227, 228, 230, 230, 230, 228, 228, 229, 230, 231, 230, 229, 230, 230, 230, 230, 229, 230, 230, 230, 231, 230, 230, 230, 230, 231, 231, 229, 230, 230, 231, 231, 230, 230, 230, 230, 230, 231, 230, 229, 230, 231, 231, 230, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 231, 230, 230, 232, 232, 232, 231, 231, 232, 232, 232, 232, 231, 231, 233, 232, 233, 232, 232, 232, 234, 234, 234, 234, 234, 235, 236, 236, 232, 227, 211, 161, 161, 157, 156, 158, 163, 159, 153, 151, 140, 144, 140, 144, 136, 150, 182, 187, 189, 166, 160, 175, 150, 82, 49, 46, 58, 79, 142, 167, 151, 59, 129, 166, 160, 98, 58, 117, 161, 166, 132, 156, 71, 42, 45, 68, 147, 146, 43, 42, 53, 135, 153, 101, 52, 52, 68, 129, 213, 231, 235, 236, 236, 234, 224, 187, 133, 54, 65, 50, 46, 56, 108, 209, 229, 229, 229, 229, 230, 231, 231, 230, 228, 229, 231, 232, 230, 230, 229, 230, 229, 230, 229, 229, 230, 231, 231, 229, 229, 228, 230, 230, 231, 229, 230, 229, 231, 231, 230, 229, 225, 222, 217, 224, 223, 219, 217, 125, 215, 224, 223, 221, 224, 220, 224, 224, 225, 226, 226, 225, 228, 227, 227, 227, 225, 228, 228, 228, 226, 227, 228, 228, 227, 227, 226, 226, 227, 228, 227, 226, 225, 227, 228, 228, 225, 226, 227, 229, 230, 230, 228, 229, 230, 231, 231, 229, 230, 229, 230, 230, 229, 229, 229, 229, 230, 230, 230, 230, 229, 231, 232, 231, 229, 230, 230, 231, 231, 230, 230, 229, 230, 230, 231, 229, 229, 229, 231, 230, 231, 230, 230, 230, 232, 231, 230, 229, 230, 231, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 230, 231, 230, 232, 231, 232, 231, 231, 231, 233, 233, 232, 232, 232, 233, 233, 233, 232, 233, 233, 234, 234, 234, 234, 234, 235, 236, 235, 231, 222, 175, 171, 165, 167, 160, 162, 162, 155, 149, 146, 139, 149, 140, 133, 137, 167, 192, 199, 185, 158, 175, 164, 105, 51, 38, 42, 50, 75, 129, 171, 157, 69, 106, 165, 158, 91, 76, 97, 167, 166, 78, 150, 105, 45, 48, 75, 146, 140, 44, 46, 56, 131, 165, 122, 42, 39, 48, 72, 120, 208, 232, 235, 236, 236, 232, 222, 181, 121, 52, 48, 47, 61, 137, 214, 227, 229, 229, 229, 230, 230, 231, 230, 229, 229, 231, 231, 230, 230, 230, 231, 231, 231, 229, 228, 229, 230, 231, 230, 228, 228, 229, 230, 231, 230, 230, 230, 231, 230, 230, 229, 224, 222, 218, 228, 223, 220, 219, 135, 213, 223, 223, 223, 224, 221, 224, 223, 225, 226, 224, 225, 225, 227, 226, 224, 224, 226, 226, 227, 227, 225, 226, 225, 226, 228, 227, 227, 227, 229, 227, 226, 227, 227, 228, 229, 228, 226, 227, 229, 230, 230, 229, 229, 229, 231, 231, 230, 229, 229, 230, 230, 229, 229, 228, 229, 229, 230, 230, 230, 229, 230, 231, 231, 229, 230, 230, 231, 231, 231, 229, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 229, 230, 230, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 232, 232, 232, 230, 231, 231, 232, 232, 232, 231, 231, 232, 233, 233, 232, 233, 233, 234, 234, 235, 234, 234, 235, 235, 233, 227, 180, 174, 169, 167, 162, 167, 165, 155, 152, 149, 146, 148, 144, 134, 134, 161, 187, 200, 198, 169, 171, 178, 133, 55, 52, 45, 46, 48, 83, 99, 177, 168, 88, 91, 166, 163, 64, 92, 88, 160, 163, 66, 91, 137, 87, 65, 101, 157, 99, 38, 39, 61, 110, 160, 126, 40, 34, 39, 47, 67, 112, 210, 232, 235, 236, 235, 231, 217, 168, 107, 50, 49, 59, 112, 189, 223, 228, 229, 229, 229, 230, 231, 230, 229, 229, 231, 231, 231, 230, 229, 230, 231, 231, 229, 228, 227, 230, 231, 230, 229, 228, 229, 230, 231, 230, 229, 229, 231, 229, 228, 230, 226, 223, 219, 228, 224, 225, 222, 119, 212, 224, 223, 223, 221, 221, 220, 224, 227, 225, 225, 226, 227, 226, 225, 224, 226, 226, 228, 228, 227, 225, 227, 228, 226, 227, 227, 227, 228, 230, 229, 228, 227, 226, 229, 228, 228, 228, 228, 229, 230, 230, 229, 230, 229, 231, 231, 230, 228, 229, 230, 230, 230, 229, 229, 229, 230, 230, 229, 229, 229, 230, 230, 231, 230, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 230, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 232, 231, 230, 230, 232, 232, 232, 231, 231, 231, 232, 232, 231, 232, 231, 232, 233, 232, 231, 232, 232, 233, 233, 233, 233, 233, 234, 234, 235, 234, 234, 235, 234, 230, 196, 176, 170, 169, 168, 166, 166, 162, 157, 149, 144, 150, 150, 130, 127, 145, 182, 193, 201, 187, 164, 185, 163, 81, 47, 46, 44, 47, 48, 60, 80, 174, 177, 87, 70, 160, 164, 68, 77, 111, 150, 156, 73, 51, 67, 82, 101, 139, 114, 48, 39, 41, 60, 97, 162, 135, 39, 34, 41, 38, 48, 72, 124, 217, 234, 235, 236, 234, 228, 209, 155, 79, 47, 50, 73, 140, 204, 224, 228, 228, 229, 231, 230, 230, 229, 230, 231, 231, 231, 229, 229, 229, 230, 231, 229, 229, 229, 229, 230, 231, 230, 228, 229, 231, 231, 231, 230, 229, 229, 230, 229, 228, 225, 223, 218, 228, 223, 224, 222, 126, 210, 221, 222, 223, 221, 223, 223, 225, 227, 224, 226, 225, 227, 226, 227, 226, 224, 226, 227, 227, 226, 227, 228, 226, 225, 226, 226, 226, 227, 229, 229, 226, 226, 228, 229, 228, 228, 228, 228, 229, 230, 229, 229, 229, 229, 230, 231, 230, 229, 229, 230, 231, 230, 229, 229, 229, 231, 230, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 232, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 231, 232, 232, 232, 233, 232, 231, 232, 233, 233, 233, 233, 233, 233, 235, 234, 235, 235, 234, 234, 231, 216, 177, 174, 173, 170, 176, 172, 171, 159, 149, 154, 152, 155, 154, 128, 136, 170, 193, 199, 201, 174, 179, 177, 119, 50, 46, 46, 44, 43, 44, 56, 68, 158, 172, 92, 62, 161, 164, 71, 64, 118, 141, 152, 82, 53, 73, 106, 97, 63, 48, 48, 41, 44, 50, 80, 158, 142, 44, 37, 38, 36, 39, 53, 72, 146, 225, 234, 236, 235, 232, 226, 194, 134, 57, 46, 56, 84, 160, 212, 226, 227, 227, 229, 231, 230, 230, 231, 231, 231, 230, 229, 229, 230, 231, 231, 230, 229, 229, 228, 230, 230, 230, 227, 230, 231, 232, 231, 229, 228, 230, 228, 228, 227, 225, 224, 219, 227, 224, 221, 222, 115, 212, 224, 221, 220, 221, 221, 225, 226, 226, 223, 227, 226, 227, 227, 226, 224, 224, 226, 228, 228, 227, 227, 228, 227, 226, 227, 228, 228, 228, 228, 229, 228, 227, 227, 229, 228, 229, 228, 228, 228, 229, 230, 229, 230, 230, 230, 231, 230, 229, 230, 230, 231, 230, 229, 229, 229, 231, 231, 230, 230, 230, 231, 231, 232, 230, 230, 230, 231, 231, 231, 229, 230, 230, 231, 230, 230, 230, 229, 231, 231, 230, 230, 230, 230, 231, 231, 230, 229, 229, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 232, 230, 230, 231, 232, 232, 231, 231, 230, 231, 232, 232, 231, 231, 231, 233, 233, 232, 231, 231, 233, 233, 233, 232, 233, 233, 235, 234, 235, 235, 233, 231, 227, 178, 183, 174, 173, 173, 175, 172, 166, 155, 155, 156, 165, 169, 160, 148, 154, 185, 200, 199, 189, 170, 186, 158, 64, 54, 43, 49, 48, 42, 48, 58, 66, 158, 170, 95, 64, 165, 165, 77, 58, 81, 155, 138, 86, 70, 117, 68, 46, 48, 41, 41, 39, 41, 51, 68, 156, 144, 63, 36, 35, 38, 35, 41, 57, 80, 180, 231, 235, 235, 234, 232, 223, 174, 105, 46, 55, 61, 108, 188, 220, 228, 227, 229, 230, 230, 230, 231, 231, 231, 230, 229, 229, 231, 230, 231, 230, 229, 229, 230, 230, 230, 230, 228, 230, 231, 230, 229, 227, 229, 230, 230, 227, 228, 223, 220, 216, 227, 222, 220, 224, 122, 214, 226, 224, 221, 222, 221, 226, 227, 226, 223, 225, 225, 226, 227, 224, 226, 224, 228, 228, 227, 228, 227, 228, 228, 229, 228, 228, 227, 229, 229, 229, 228, 226, 228, 230, 229, 228, 228, 226, 227, 229, 229, 230, 229, 229, 230, 230, 230, 229, 229, 231, 230, 230, 229, 228, 229, 231, 231, 230, 230, 230, 231, 230, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 232, 231, 230, 230, 232, 232, 232, 231, 231, 231, 233, 233, 232, 231, 231, 232, 233, 233, 233, 233, 233, 234, 234, 235, 234, 232, 229, 195, 181, 179, 177, 174, 176, 176, 167, 161, 158, 158, 170, 170, 170, 178, 161, 173, 194, 199, 199, 173, 178, 178, 113, 48, 47, 49, 47, 52, 43, 46, 56, 61, 162, 174, 89, 74, 156, 164, 77, 56, 64, 155, 130, 88, 136, 145, 132, 106, 103, 89, 95, 52, 45, 48, 62, 159, 148, 58, 39, 39, 38, 38, 40, 56, 61, 88, 200, 233, 235, 235, 235, 229, 209, 148, 64, 46, 52, 72, 141, 203, 221, 226, 228, 230, 230, 230, 231, 231, 230, 230, 229, 229, 230, 230, 231, 230, 230, 230, 230, 231, 229, 229, 229, 230, 231, 230, 230, 229, 228, 229, 229, 229, 228, 224, 222, 215, 229, 223, 220, 224, 124, 216, 226, 226, 223, 222, 223, 225, 228, 226, 225, 227, 227, 224, 227, 225, 226, 227, 228, 230, 228, 228, 227, 226, 228, 227, 228, 228, 228, 229, 228, 228, 229, 228, 228, 230, 229, 227, 228, 228, 227, 229, 229, 230, 229, 229, 230, 231, 229, 229, 229, 230, 231, 229, 229, 229, 229, 231, 231, 230, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 229, 230, 231, 231, 231, 229, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 229, 229, 230, 230, 230, 231, 229, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 232, 230, 230, 230, 232, 232, 232, 231, 231, 232, 233, 233, 232, 232, 232, 233, 234, 233, 232, 233, 233, 234, 235, 235, 233, 229, 221, 173, 179, 178, 176, 181, 181, 179, 169, 162, 158, 167, 174, 179, 176, 175, 181, 188, 196, 202, 191, 167, 183, 165, 70, 50, 51, 57, 46, 45, 41, 42, 51, 54, 147, 168, 105, 63, 156, 162, 87, 56, 59, 149, 147, 112, 132, 166, 174, 165, 162, 166, 151, 55, 43, 50, 58, 162, 154, 63, 35, 37, 34, 36, 40, 38, 46, 67, 121, 221, 235, 235, 236, 233, 225, 184, 115, 50, 47, 58, 88, 170, 212, 224, 227, 230, 230, 230, 230, 232, 230, 230, 229, 230, 230, 231, 231, 229, 230, 230, 231, 230, 229, 229, 229, 230, 231, 230, 229, 230, 229, 230, 230, 231, 229, 225, 222, 214, 226, 222, 221, 226, 125, 218, 225, 226, 222, 222, 224, 226, 227, 228, 226, 226, 226, 226, 227, 226, 226, 228, 228, 230, 228, 228, 227, 227, 227, 227, 226, 227, 228, 230, 229, 229, 228, 228, 229, 229, 230, 229, 229, 227, 228, 230, 230, 229, 230, 229, 230, 231, 229, 229, 229, 230, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 230, 231, 230, 230, 229, 231, 231, 231, 229, 230, 230, 231, 232, 230, 230, 230, 230, 231, 231, 230, 229, 229, 231, 231, 231, 230, 230, 230, 231, 232, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 231, 231, 230, 230, 232, 231, 232, 231, 231, 232, 233, 233, 232, 232, 232, 233, 233, 234, 233, 233, 233, 235, 236, 234, 232, 229, 186, 180, 180, 179, 174, 175, 178, 172, 168, 162, 159, 172, 176, 179, 178, 180, 181, 187, 198, 203, 180, 176, 177, 140, 85, 80, 130, 131, 62, 43, 47, 42, 51, 55, 144, 172, 113, 59, 153, 173, 104, 54, 55, 142, 125, 97, 101, 128, 141, 143, 149, 142, 100, 49, 41, 50, 58, 152, 160, 58, 36, 39, 41, 43, 47, 41, 46, 59, 85, 173, 230, 235, 236, 236, 230, 212, 155, 73, 45, 49, 67, 123, 189, 219, 225, 230, 230, 230, 230, 231, 230, 229, 229, 229, 230, 230, 230, 230, 229, 230, 231, 231, 230, 229, 229, 230, 231, 230, 228, 229, 228, 229, 229, 229, 230, 225, 223, 218, 225, 222, 220, 224, 114, 217, 225, 227, 224, 223, 225, 227, 227, 226, 226, 227, 226, 227, 228, 228, 226, 228, 228, 229, 228, 229, 227, 228, 228, 227, 227, 227, 227, 230, 229, 229, 228, 229, 229, 230, 230, 229, 229, 228, 228, 230, 230, 229, 230, 230, 231, 231, 230, 229, 229, 230, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 229, 229, 229, 231, 231, 231, 229, 230, 230, 232, 232, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 230, 230, 232, 232, 232, 231, 231, 232, 233, 233, 232, 232, 232, 233, 233, 233, 232, 233, 234, 235, 235, 233, 229, 218, 172, 180, 180, 176, 171, 180, 175, 171, 165, 157, 167, 179, 180, 182, 179, 178, 182, 193, 201, 195, 174, 184, 180, 104, 170, 103, 169, 168, 75, 48, 48, 42, 52, 55, 141, 170, 131, 62, 140, 180, 134, 54, 57, 90, 56, 54, 71, 81, 57, 53, 64, 78, 46, 38, 37, 50, 52, 153, 165, 67, 42, 60, 126, 94, 90, 115, 70, 54, 83, 125, 212, 234, 236, 236, 234, 226, 182, 126, 51, 49, 57, 80, 160, 213, 225, 229, 230, 230, 230, 230, 230, 230, 229, 229, 229, 230, 231, 229, 228, 230, 229, 230, 230, 228, 228, 229, 231, 228, 229, 229, 229, 230, 230, 229, 229, 226, 225, 221, 228, 222, 222, 223, 114, 218, 227, 226, 223, 225, 226, 225, 227, 228, 225, 228, 227, 229, 227, 228, 228, 229, 229, 229, 229, 228, 227, 229, 230, 228, 228, 227, 228, 230, 229, 229, 229, 229, 230, 230, 230, 229, 228, 229, 229, 230, 231, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 231, 230, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 230, 230, 229, 230, 231, 231, 230, 230, 229, 231, 232, 231, 230, 230, 230, 232, 232, 231, 230, 230, 231, 232, 232, 231, 230, 230, 232, 233, 232, 231, 232, 232, 232, 233, 232, 232, 232, 233, 233, 233, 232, 233, 234, 236, 234, 232, 227, 184, 174, 179, 178, 177, 175, 179, 175, 172, 161, 163, 178, 180, 180, 180, 184, 184, 190, 199, 202, 196, 167, 186, 159, 71, 88, 103, 161, 170, 83, 48, 77, 68, 66, 57, 112, 137, 111, 56, 113, 152, 125, 54, 66, 100, 48, 48, 68, 91, 93, 50, 51, 82, 60, 41, 45, 67, 67, 136, 158, 73, 46, 118, 139, 48, 51, 105, 151, 77, 98, 192, 158, 230, 235, 236, 236, 229, 213, 159, 76, 49, 52, 63, 119, 196, 223, 229, 229, 230, 229, 230, 231, 230, 229, 228, 229, 230, 230, 229, 228, 229, 230, 230, 229, 229, 229, 231, 230, 231, 230, 230, 229, 230, 230, 230, 228, 226, 226, 220, 229, 223, 220, 222, 129, 216, 228, 228, 225, 225, 228, 227, 226, 225, 226, 226, 227, 230, 227, 228, 228, 228, 229, 229, 228, 227, 226, 229, 229, 229, 229, 228, 228, 229, 229, 229, 229, 229, 229, 231, 231, 230, 228, 229, 229, 230, 230, 229, 230, 229, 230, 230, 229, 230, 230, 231, 231, 231, 230, 230, 230, 231, 230, 230, 229, 229, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 230, 229, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 230, 232, 232, 230, 230, 230, 232, 231, 231, 231, 230, 231, 232, 232, 231, 231, 230, 231, 232, 232, 232, 232, 232, 233, 233, 233, 232, 232, 233, 234, 233, 233, 233, 234, 235, 233, 229, 223, 164, 177, 180, 181, 173, 179, 175, 169, 171, 165, 173, 180, 182, 181, 182, 184, 188, 189, 202, 206, 191, 177, 182, 149, 63, 59, 90, 160, 174, 99, 108, 128, 58, 120, 92, 57, 47, 51, 48, 46, 54, 55, 58, 90, 135, 52, 50, 100, 98, 96, 71, 63, 131, 122, 39, 44, 60, 70, 54, 61, 46, 46, 144, 131, 46, 50, 72, 151, 117, 57, 87, 97, 208, 235, 236, 236, 232, 225, 186, 115, 50, 47, 57, 85, 172, 219, 229, 230, 229, 230, 231, 231, 230, 229, 229, 230, 230, 230, 229, 229, 230, 230, 231, 229, 230, 229, 230, 231, 231, 230, 229, 230, 230, 230, 229, 228, 225, 224, 222, 225, 222, 217, 221, 121, 216, 226, 226, 225, 226, 226, 228, 226, 226, 226, 227, 228, 229, 229, 228, 228, 227, 229, 228, 228, 228, 228, 229, 229, 229, 229, 229, 227, 229, 229, 229, 229, 229, 229, 230, 231, 229, 229, 229, 229, 230, 231, 230, 229, 230, 230, 230, 230, 230, 229, 230, 230, 230, 230, 230, 229, 231, 231, 230, 229, 229, 231, 230, 230, 229, 229, 230, 231, 231, 231, 230, 229, 230, 231, 230, 230, 229, 230, 231, 231, 230, 229, 229, 230, 231, 230, 229, 229, 229, 230, 231, 230, 230, 230, 230, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 232, 233, 233, 232, 232, 232, 232, 234, 233, 233, 233, 234, 235, 233, 228, 201, 178, 175, 183, 180, 176, 176, 174, 169, 173, 168, 178, 184, 183, 186, 186, 185, 187, 193, 205, 207, 182, 180, 176, 121, 53, 59, 59, 152, 182, 108, 153, 120, 61, 101, 152, 63, 47, 47, 45, 42, 42, 48, 49, 51, 94, 50, 47, 51, 58, 54, 61, 82, 75, 62, 42, 45, 46, 48, 99, 93, 43, 42, 137, 143, 48, 51, 73, 142, 135, 46, 59, 83, 161, 232, 236, 237, 234, 228, 209, 150, 61, 48, 50, 69, 137, 207, 227, 229, 230, 230, 231, 231, 230, 230, 230, 230, 231, 230, 229, 229, 230, 230, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 230, 230, 228, 230, 225, 225, 221, 228, 222, 219, 223, 123, 218, 226, 226, 224, 226, 226, 228, 227, 226, 226, 226, 227, 229, 229, 228, 228, 227, 228, 228, 229, 229, 228, 230, 230, 229, 229, 228, 229, 230, 230, 230, 229, 229, 229, 230, 230, 230, 230, 230, 230, 230, 231, 230, 230, 230, 230, 231, 230, 230, 229, 231, 231, 230, 230, 230, 230, 231, 231, 229, 228, 229, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 229, 230, 231, 231, 231, 230, 230, 229, 230, 231, 230, 230, 230, 230, 231, 231, 229, 229, 230, 231, 231, 231, 230, 230, 231, 232, 231, 231, 231, 231, 232, 232, 232, 232, 232, 232, 233, 233, 232, 232, 232, 233, 234, 234, 233, 234, 235, 234, 232, 229, 175, 177, 176, 182, 178, 179, 178, 173, 175, 172, 171, 178, 181, 186, 186, 187, 187, 188, 200, 207, 205, 180, 190, 172, 110, 53, 53, 59, 141, 182, 123, 164, 112, 66, 84, 162, 99, 51, 46, 46, 39, 43, 44, 48, 57, 109, 110, 49, 48, 43, 47, 52, 57, 138, 78, 41, 42, 43, 38, 38, 39, 41, 48, 96, 150, 91, 62, 72, 148, 110, 49, 51, 76, 106, 218, 236, 236, 235, 230, 222, 178, 82, 48, 44, 63, 95, 192, 224, 229, 230, 230, 231, 231, 230, 230, 229, 230, 230, 231, 229, 230, 230, 230, 230, 230, 230, 229, 230, 231, 230, 230, 229, 229, 231, 230, 229, 229, 226, 225, 218, 229, 224, 223, 223, 125, 217, 225, 226, 224, 226, 226, 228, 228, 227, 227, 227, 228, 229, 229, 229, 229, 228, 229, 228, 229, 228, 227, 229, 230, 230, 230, 229, 230, 230, 230, 230, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 229, 229, 231, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 229, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 230, 231, 231, 232, 232, 232, 231, 232, 232, 233, 232, 232, 231, 233, 234, 234, 233, 234, 234, 233, 229, 218, 171, 178, 178, 182, 178, 178, 178, 174, 175, 177, 179, 180, 187, 183, 190, 189, 189, 196, 205, 203, 206, 182, 184, 167, 79, 48, 53, 57, 136, 184, 137, 166, 122, 63, 70, 162, 124, 50, 43, 43, 43, 45, 50, 51, 47, 89, 93, 59, 50, 51, 53, 59, 67, 121, 104, 57, 45, 41, 41, 39, 39, 43, 46, 51, 95, 123, 96, 109, 124, 56, 48, 50, 66, 84, 183, 234, 236, 235, 233, 227, 200, 122, 49, 44, 52, 78, 168, 219, 229, 230, 230, 230, 231, 230, 230, 230, 230, 230, 230, 229, 230, 230, 231, 231, 231, 230, 229, 230, 230, 230, 230, 230, 229, 229, 230, 230, 230, 227, 225, 221, 229, 225, 223, 224, 129, 219, 226, 227, 224, 224, 225, 226, 225, 226, 226, 228, 228, 230, 230, 229, 228, 227, 228, 230, 229, 229, 228, 229, 231, 230, 230, 230, 229, 230, 230, 230, 229, 230, 230, 232, 231, 230, 230, 229, 231, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 230, 230, 230, 229, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 229, 229, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 231, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 233, 231, 231, 231, 232, 233, 233, 231, 232, 233, 234, 234, 233, 234, 233, 233, 229, 193, 177, 178, 182, 182, 180, 183, 185, 177, 178, 175, 180, 182, 188, 187, 188, 193, 192, 196, 204, 207, 205, 178, 186, 159, 59, 52, 52, 60, 124, 183, 145, 155, 139, 62, 66, 151, 129, 52, 49, 45, 45, 45, 43, 43, 49, 48, 78, 128, 79, 61, 72, 84, 110, 69, 55, 64, 62, 48, 41, 42, 45, 40, 44, 46, 50, 77, 102, 85, 54, 50, 48, 48, 61, 81, 132, 229, 235, 235, 234, 228, 216, 151, 57, 44, 48, 68, 132, 207, 228, 229, 230, 231, 231, 230, 230, 229, 230, 230, 230, 230, 230, 230, 231, 231, 230, 230, 230, 230, 230, 231, 229, 230, 229, 228, 229, 230, 230, 228, 227, 221, 226, 224, 223, 224, 140, 219, 228, 225, 226, 225, 227, 226, 227, 227, 227, 228, 227, 229, 230, 229, 227, 227, 229, 230, 229, 228, 229, 229, 230, 230, 230, 229, 228, 231, 230, 230, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 230, 230, 229, 229, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 229, 230, 229, 231, 231, 231, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 232, 231, 231, 231, 232, 232, 233, 232, 231, 232, 232, 233, 233, 232, 232, 233, 234, 234, 233, 234, 233, 232, 229, 179, 178, 175, 186, 181, 178, 186, 182, 175, 178, 181, 182, 184, 183, 189, 189, 193, 195, 197, 207, 209, 200, 181, 187, 148, 55, 50, 51, 61, 122, 177, 149, 134, 152, 65, 67, 159, 100, 48, 46, 41, 40, 41, 42, 46, 43, 49, 48, 102, 90, 128, 130, 83, 91, 46, 50, 49, 60, 57, 49, 40, 40, 44, 42, 48, 95, 87, 62, 57, 56, 67, 52, 49, 57, 74, 104, 216, 235, 235, 235, 231, 224, 176, 82, 44, 45, 75, 94, 191, 224, 229, 230, 230, 231, 230, 229, 229, 230, 230, 230, 230, 229, 230, 231, 231, 231, 229, 229, 230, 231, 231, 229, 229, 229, 229, 230, 230, 229, 227, 226, 220, 225, 222, 222, 224, 135, 220, 228, 228, 226, 225, 226, 224, 226, 227, 228, 227, 229, 229, 230, 227, 229, 228, 228, 229, 228, 229, 229, 228, 229, 230, 230, 229, 229, 231, 231, 230, 229, 230, 230, 231, 231, 230, 230, 229, 230, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 232, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 232, 231, 231, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 232, 231, 231, 231, 231, 232, 232, 232, 231, 232, 233, 233, 232, 232, 232, 234, 234, 234, 234, 233, 233, 229, 220, 168, 175, 179, 188, 177, 188, 185, 182, 180, 179, 183, 185, 184, 181, 187, 189, 194, 196, 202, 206, 210, 201, 181, 181, 137, 48, 49, 52, 64, 106, 176, 159, 74, 152, 91, 84, 146, 59, 41, 44, 41, 42, 39, 41, 41, 46, 47, 50, 51, 93, 78, 67, 71, 61, 51, 45, 42, 51, 43, 56, 46, 37, 49, 46, 64, 158, 162, 161, 155, 153, 123, 50, 55, 58, 72, 95, 188, 234, 235, 235, 233, 227, 191, 111, 50, 48, 56, 83, 176, 222, 230, 230, 231, 231, 231, 229, 230, 229, 231, 231, 229, 229, 230, 231, 230, 230, 230, 230, 230, 228, 230, 229, 229, 227, 230, 230, 231, 229, 228, 225, 222, 226, 224, 224, 224, 144, 219, 228, 227, 226, 226, 226, 227, 228, 228, 229, 229, 229, 230, 230, 228, 227, 227, 228, 230, 228, 228, 228, 228, 229, 230, 229, 229, 229, 231, 231, 230, 229, 229, 230, 231, 231, 230, 230, 229, 232, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 230, 229, 230, 231, 231, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 231, 230, 230, 230, 231, 231, 231, 229, 230, 231, 232, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 231, 231, 231, 231, 231, 233, 232, 231, 231, 232, 233, 233, 233, 232, 232, 233, 234, 234, 234, 233, 232, 228, 208, 175, 180, 180, 187, 181, 184, 187, 182, 184, 184, 184, 187, 184, 184, 193, 189, 195, 192, 202, 209, 214, 199, 186, 187, 138, 52, 48, 55, 58, 74, 125, 111, 56, 67, 87, 89, 67, 47, 43, 43, 37, 45, 39, 40, 39, 36, 44, 56, 92, 179, 161, 157, 174, 159, 99, 43, 47, 45, 41, 45, 54, 49, 46, 55, 80, 154, 163, 157, 157, 144, 87, 56, 55, 62, 69, 90, 148, 232, 235, 236, 234, 228, 203, 136, 52, 50, 56, 73, 145, 215, 228, 229, 231, 230, 230, 229, 229, 229, 230, 230, 229, 230, 228, 230, 231, 230, 230, 229, 229, 230, 230, 228, 227, 229, 231, 229, 229, 228, 228, 226, 220, 228, 221, 220, 223, 130, 218, 228, 227, 224, 226, 226, 227, 229, 228, 228, 229, 230, 230, 230, 228, 227, 227, 229, 230, 229, 228, 229, 229, 230, 230, 229, 229, 229, 230, 231, 230, 228, 229, 230, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 229, 229, 230, 230, 231, 231, 229, 230, 229, 231, 231, 230, 230, 229, 231, 231, 231, 229, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 232, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 232, 230, 230, 231, 232, 233, 232, 231, 231, 232, 233, 233, 233, 232, 232, 234, 234, 234, 234, 233, 232, 230, 191, 178, 179, 184, 186, 185, 187, 187, 182, 180, 180, 187, 184, 188, 189, 196, 192, 192, 193, 203, 210, 211, 199, 196, 189, 138, 55, 49, 49, 54, 50, 54, 52, 47, 51, 45, 47, 40, 40, 39, 41, 41, 56, 40, 40, 37, 40, 50, 56, 169, 170, 176, 180, 179, 150, 108, 49, 55, 52, 46, 53, 53, 53, 61, 53, 51, 61, 66, 56, 59, 57, 49, 55, 56, 61, 68, 90, 120, 223, 235, 235, 235, 229, 208, 150, 56, 52, 54, 68, 116, 206, 228, 229, 231, 231, 230, 229, 229, 230, 230, 229, 228, 229, 230, 231, 231, 231, 230, 229, 229, 230, 230, 229, 228, 229, 231, 231, 230, 229, 225, 225, 217, 228, 224, 221, 223, 146, 222, 227, 227, 226, 226, 226, 227, 227, 227, 226, 227, 229, 230, 230, 228, 228, 229, 229, 230, 229, 228, 229, 230, 230, 230, 230, 229, 230, 230, 231, 230, 229, 229, 230, 231, 231, 229, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 231, 232, 232, 230, 231, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 233, 232, 231, 231, 232, 233, 233, 232, 232, 232, 234, 234, 234, 234, 233, 231, 230, 189, 183, 183, 184, 188, 182, 191, 185, 177, 176, 182, 186, 191, 189, 188, 196, 192, 192, 193, 199, 208, 210, 196, 189, 185, 133, 46, 48, 53, 64, 89, 92, 89, 65, 49, 45, 44, 44, 43, 44, 39, 39, 38, 41, 39, 35, 41, 47, 61, 148, 166, 152, 137, 130, 100, 98, 52, 47, 50, 45, 47, 46, 53, 57, 63, 67, 49, 53, 47, 54, 50, 61, 64, 64, 66, 69, 84, 100, 212, 234, 235, 235, 230, 217, 159, 69, 51, 59, 69, 103, 199, 225, 229, 231, 231, 230, 230, 229, 230, 230, 231, 229, 230, 230, 231, 232, 231, 230, 229, 228, 230, 230, 229, 229, 230, 231, 231, 231, 230, 228, 225, 217, 228, 225, 220, 223, 127, 220, 228, 227, 227, 227, 228, 228, 229, 229, 228, 228, 228, 230, 230, 229, 229, 230, 230, 229, 228, 228, 229, 229, 230, 230, 230, 229, 230, 231, 231, 230, 229, 229, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 229, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 229, 229, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 233, 232, 231, 232, 232, 233, 233, 232, 232, 232, 233, 234, 234, 233, 233, 230, 230, 183, 180, 180, 186, 186, 185, 188, 183, 179, 179, 179, 186, 186, 188, 186, 192, 193, 190, 196, 202, 210, 211, 196, 189, 189, 135, 52, 53, 70, 142, 125, 89, 123, 146, 90, 51, 40, 40, 45, 43, 44, 39, 38, 44, 41, 41, 40, 48, 52, 124, 133, 126, 139, 169, 159, 131, 57, 47, 49, 46, 61, 48, 51, 47, 58, 59, 72, 67, 58, 60, 114, 142, 149, 143, 107, 68, 81, 104, 191, 233, 235, 235, 231, 221, 168, 82, 50, 52, 65, 96, 186, 224, 229, 231, 231, 230, 230, 229, 231, 230, 231, 230, 230, 230, 231, 230, 231, 229, 228, 230, 230, 230, 229, 229, 230, 231, 231, 231, 228, 228, 226, 219, 228, 224, 222, 224, 123, 217, 227, 228, 227, 227, 228, 227, 228, 229, 228, 226, 229, 230, 231, 228, 227, 228, 229, 229, 229, 228, 229, 229, 230, 230, 230, 229, 229, 231, 230, 231, 230, 229, 229, 231, 230, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 230, 231, 230, 229, 230, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 230, 230, 231, 231, 231, 231, 230, 230, 231, 232, 232, 231, 230, 231, 232, 232, 232, 231, 231, 232, 233, 232, 232, 232, 232, 233, 234, 234, 233, 233, 230, 230, 181, 181, 179, 185, 185, 184, 189, 184, 177, 179, 179, 186, 185, 185, 190, 185, 194, 192, 189, 198, 209, 211, 195, 191, 188, 142, 55, 59, 126, 165, 70, 57, 87, 140, 159, 61, 47, 46, 42, 43, 45, 38, 39, 43, 42, 44, 37, 44, 49, 54, 60, 101, 162, 173, 178, 159, 115, 56, 55, 50, 56, 56, 60, 55, 60, 65, 69, 110, 118, 81, 146, 163, 148, 163, 111, 106, 113, 127, 178, 231, 234, 234, 231, 224, 176, 90, 56, 56, 65, 90, 173, 222, 230, 231, 231, 231, 230, 230, 230, 229, 231, 230, 229, 230, 232, 231, 231, 229, 229, 230, 230, 230, 229, 229, 230, 231, 231, 230, 229, 228, 227, 219, 226, 224, 223, 223, 129, 219, 226, 227, 227, 227, 228, 229, 229, 228, 227, 228, 229, 229, 229, 226, 228, 227, 228, 229, 230, 228, 229, 230, 231, 231, 230, 229, 228, 230, 231, 230, 230, 229, 230, 231, 230, 230, 229, 229, 231, 231, 231, 229, 229, 230, 231, 231, 230, 229, 229, 230, 231, 230, 229, 230, 230, 230, 230, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 230, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 229, 230, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 232, 231, 230, 231, 232, 232, 232, 231, 231, 231, 233, 233, 232, 232, 233, 233, 234, 234, 232, 232, 230, 229, 179, 183, 182, 186, 186, 191, 190, 184, 180, 178, 179, 184, 183, 185, 187, 187, 188, 185, 188, 200, 206, 209, 199, 187, 188, 143, 56, 54, 141, 159, 59, 56, 65, 107, 166, 117, 43, 40, 39, 37, 40, 39, 37, 38, 40, 38, 40, 38, 44, 48, 57, 142, 166, 164, 163, 170, 161, 140, 143, 140, 142, 144, 148, 148, 143, 152, 153, 163, 174, 156, 150, 168, 194, 205, 200, 201, 204, 207, 210, 216, 231, 234, 232, 227, 180, 112, 57, 58, 66, 88, 166, 218, 229, 231, 231, 230, 230, 228, 230, 230, 230, 230, 230, 230, 232, 231, 230, 230, 229, 229, 228, 230, 227, 228, 229, 230, 231, 230, 230, 227, 226, 218, 227, 223, 221, 224, 118, 218, 227, 226, 225, 227, 228, 228, 228, 228, 227, 228, 228, 229, 229, 228, 228, 227, 229, 229, 229, 229, 229, 230, 230, 231, 230, 229, 228, 230, 231, 230, 229, 229, 229, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 229, 229, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 231, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 232, 232, 231, 230, 231, 231, 232, 232, 231, 232, 231, 233, 233, 233, 232, 232, 233, 234, 234, 233, 232, 230, 230, 185, 181, 182, 187, 186, 189, 192, 183, 179, 178, 179, 185, 187, 184, 183, 183, 189, 190, 188, 201, 207, 211, 203, 182, 191, 155, 61, 54, 126, 155, 72, 53, 58, 86, 161, 154, 51, 38, 40, 40, 40, 42, 41, 33, 37, 35, 39, 38, 45, 70, 68, 145, 165, 166, 140, 174, 170, 171, 169, 166, 167, 158, 158, 152, 150, 151, 146, 144, 145, 146, 128, 143, 160, 160, 168, 146, 134, 148, 158, 222, 232, 234, 233, 228, 182, 122, 59, 55, 66, 88, 154, 217, 229, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 231, 231, 230, 231, 229, 229, 230, 228, 228, 229, 228, 228, 230, 230, 230, 229, 229, 226, 220, 228, 224, 222, 224, 112, 215, 226, 218, 227, 227, 227, 228, 228, 229, 228, 228, 229, 229, 228, 227, 228, 227, 230, 229, 229, 229, 227, 229, 229, 231, 230, 229, 229, 230, 230, 230, 229, 230, 229, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 229, 230, 230, 231, 230, 229, 229, 231, 231, 231, 230, 230, 230, 232, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 231, 231, 232, 233, 232, 231, 232, 233, 233, 232, 232, 232, 233, 234, 234, 234, 232, 230, 230, 186, 183, 185, 188, 181, 186, 193, 181, 183, 179, 179, 181, 182, 182, 185, 186, 189, 189, 191, 197, 209, 217, 208, 189, 197, 166, 78, 54, 78, 152, 118, 61, 61, 76, 160, 161, 51, 43, 43, 40, 40, 42, 37, 45, 42, 39, 39, 37, 47, 53, 59, 150, 174, 176, 163, 169, 163, 120, 99, 93, 90, 85, 79, 67, 68, 62, 61, 59, 63, 83, 101, 110, 96, 92, 140, 144, 90, 144, 168, 225, 234, 234, 232, 226, 185, 119, 61, 61, 68, 100, 147, 215, 228, 230, 231, 230, 229, 229, 230, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 229, 229, 230, 229, 229, 228, 230, 230, 230, 230, 230, 226, 220, 227, 224, 224, 223, 146, 217, 227, 224, 225, 225, 225, 227, 228, 230, 227, 228, 228, 229, 227, 228, 228, 228, 229, 230, 230, 229, 228, 228, 230, 230, 231, 230, 230, 230, 231, 230, 229, 229, 229, 231, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 231, 230, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 232, 230, 231, 232, 232, 233, 232, 232, 231, 233, 233, 233, 232, 232, 233, 234, 234, 234, 232, 231, 230, 185, 182, 184, 186, 182, 184, 186, 182, 182, 182, 180, 183, 184, 184, 187, 186, 187, 190, 194, 199, 212, 218, 213, 187, 195, 168, 68, 44, 55, 86, 124, 96, 76, 63, 159, 156, 51, 42, 42, 44, 43, 43, 43, 41, 41, 41, 41, 39, 44, 49, 59, 96, 161, 170, 170, 166, 134, 59, 50, 48, 49, 54, 56, 51, 52, 50, 52, 55, 57, 105, 94, 57, 67, 72, 99, 137, 95, 98, 115, 222, 233, 234, 232, 227, 189, 124, 63, 57, 69, 95, 148, 211, 229, 231, 231, 231, 230, 229, 230, 230, 230, 230, 230, 230, 231, 231, 231, 229, 229, 228, 229, 230, 229, 228, 228, 229, 230, 230, 229, 229, 226, 220, 226, 225, 224, 224, 134, 216, 228, 227, 225, 225, 227, 227, 229, 230, 227, 227, 227, 228, 229, 226, 227, 226, 229, 230, 230, 228, 229, 228, 230, 231, 231, 230, 229, 230, 231, 231, 230, 229, 229, 231, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 231, 230, 230, 229, 230, 230, 231, 231, 230, 230, 229, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 231, 229, 230, 231, 231, 231, 230, 230, 230, 231, 232, 230, 230, 230, 231, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 232, 232, 233, 233, 233, 232, 232, 234, 235, 234, 234, 233, 231, 230, 185, 177, 179, 189, 181, 182, 193, 182, 179, 179, 183, 182, 184, 184, 187, 188, 185, 190, 194, 200, 211, 222, 216, 192, 199, 179, 90, 49, 54, 103, 113, 58, 58, 79, 163, 111, 43, 39, 44, 43, 43, 43, 42, 57, 42, 39, 40, 40, 47, 56, 68, 57, 106, 146, 157, 156, 74, 54, 49, 49, 48, 49, 51, 48, 49, 50, 53, 55, 59, 96, 95, 55, 57, 67, 107, 158, 112, 120, 119, 220, 233, 234, 232, 224, 179, 119, 58, 66, 68, 97, 152, 217, 229, 231, 231, 230, 230, 229, 230, 231, 230, 231, 229, 230, 231, 231, 231, 230, 230, 229, 230, 230, 229, 228, 228, 229, 230, 231, 229, 229, 226, 220, 227, 224, 223, 225, 125, 217, 226, 225, 224, 225, 226, 226, 227, 229, 226, 226, 226, 228, 228, 226, 226, 227, 229, 230, 230, 229, 228, 229, 230, 231, 230, 229, 230, 230, 230, 230, 230, 229, 230, 230, 231, 231, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 229, 230, 230, 232, 231, 230, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 229, 229, 231, 230, 231, 230, 230, 230, 231, 230, 229, 229, 229, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 232, 233, 233, 233, 232, 232, 234, 234, 234, 233, 233, 231, 230, 195, 178, 181, 186, 185, 187, 192, 184, 178, 178, 177, 182, 184, 184, 186, 186, 192, 194, 194, 204, 212, 222, 216, 194, 196, 183, 100, 50, 52, 112, 148, 79, 64, 134, 144, 55, 45, 45, 43, 42, 38, 41, 43, 45, 45, 44, 41, 40, 44, 46, 47, 46, 59, 70, 128, 158, 106, 54, 43, 51, 50, 50, 49, 45, 51, 52, 54, 54, 58, 65, 108, 75, 61, 71, 138, 146, 76, 99, 122, 204, 230, 233, 231, 224, 179, 116, 61, 63, 77, 108, 156, 217, 229, 231, 232, 231, 229, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 230, 229, 228, 229, 230, 230, 230, 230, 226, 229, 225, 220, 227, 225, 223, 224, 130, 220, 224, 226, 224, 224, 225, 226, 227, 228, 226, 226, 227, 228, 228, 227, 228, 228, 227, 230, 228, 228, 228, 229, 230, 231, 229, 229, 230, 231, 230, 231, 230, 229, 229, 230, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 229, 230, 230, 232, 231, 231, 229, 229, 230, 230, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 232, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 231, 232, 230, 234, 231, 231, 231, 230, 231, 231, 231, 231, 230, 230, 232, 232, 231, 230, 230, 231, 231, 231, 231, 230, 231, 232, 232, 231, 231, 231, 232, 233, 233, 233, 232, 232, 233, 234, 234, 233, 233, 231, 230, 191, 179, 181, 189, 187, 185, 191, 185, 181, 179, 181, 182, 181, 189, 187, 189, 192, 194, 196, 202, 210, 221, 222, 197, 196, 204, 127, 49, 47, 53, 99, 110, 110, 118, 57, 43, 44, 41, 39, 40, 40, 40, 43, 44, 47, 40, 46, 39, 41, 47, 42, 47, 50, 63, 88, 163, 147, 58, 50, 47, 51, 47, 49, 49, 46, 50, 49, 58, 56, 60, 69, 103, 96, 111, 124, 82, 74, 86, 112, 221, 232, 230, 227, 217, 175, 111, 67, 65, 79, 116, 163, 217, 230, 230, 231, 231, 230, 229, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 230, 229, 230, 230, 228, 229, 229, 230, 228, 228, 227, 225, 219, 226, 223, 221, 225, 124, 220, 225, 228, 225, 225, 226, 227, 229, 229, 226, 225, 227, 228, 228, 227, 227, 227, 228, 230, 230, 229, 229, 230, 230, 230, 229, 229, 229, 231, 231, 230, 229, 229, 229, 230, 230, 229, 228, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 229, 230, 230, 231, 230, 230, 230, 231, 231, 230, 230, 229, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 232, 231, 230, 230, 232, 232, 231, 230, 230, 230, 231, 230, 231, 230, 230, 231, 232, 231, 230, 230, 230, 232, 232, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 231, 231, 231, 231, 231, 232, 232, 231, 231, 232, 233, 233, 232, 232, 233, 232, 234, 234, 233, 233, 232, 231, 203, 184, 184, 192, 191, 188, 192, 186, 182, 179, 179, 183, 187, 185, 188, 190, 193, 192, 193, 200, 212, 218, 224, 205, 194, 220, 164, 53, 46, 45, 47, 49, 47, 46, 43, 41, 42, 48, 41, 47, 42, 41, 43, 40, 46, 43, 42, 43, 40, 41, 45, 58, 48, 92, 66, 138, 161, 105, 49, 58, 52, 49, 48, 49, 53, 51, 51, 53, 50, 50, 53, 61, 58, 62, 63, 58, 69, 94, 117, 224, 234, 233, 229, 217, 172, 109, 67, 68, 83, 122, 164, 218, 230, 231, 231, 231, 230, 230, 231, 231, 230, 230, 230, 230, 232, 231, 230, 230, 229, 230, 230, 230, 230, 226, 228, 230, 231, 229, 228, 227, 226, 221, 223, 221, 221, 225, 135, 217, 226, 226, 226, 224, 226, 226, 228, 228, 226, 227, 227, 229, 230, 227, 229, 230, 229, 230, 230, 228, 229, 229, 231, 230, 229, 229, 229, 230, 230, 231, 229, 229, 229, 231, 231, 229, 229, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 230, 230, 231, 230, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 230, 231, 230, 230, 231, 232, 232, 231, 230, 231, 232, 232, 231, 230, 229, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 232, 233, 233, 232, 232, 232, 233, 234, 234, 234, 233, 233, 232, 209, 186, 185, 188, 189, 186, 188, 188, 183, 180, 184, 184, 189, 182, 186, 186, 193, 186, 194, 198, 204, 213, 223, 212, 191, 224, 191, 69, 43, 38, 41, 41, 46, 55, 67, 58, 47, 44, 40, 46, 40, 39, 43, 40, 40, 40, 41, 40, 43, 45, 50, 79, 49, 96, 64, 114, 160, 142, 54, 53, 48, 51, 50, 51, 51, 53, 52, 49, 54, 55, 76, 88, 66, 52, 56, 57, 71, 85, 130, 227, 234, 233, 229, 214, 163, 102, 71, 72, 88, 118, 167, 222, 230, 231, 229, 230, 229, 230, 231, 230, 231, 230, 230, 230, 232, 231, 231, 229, 230, 230, 231, 231, 229, 228, 229, 230, 230, 229, 226, 228, 224, 222, 224, 222, 219, 224, 132, 219, 227, 227, 227, 225, 225, 226, 228, 228, 226, 226, 228, 228, 229, 228, 228, 228, 229, 230, 230, 229, 228, 229, 230, 229, 229, 228, 230, 230, 230, 230, 229, 229, 229, 231, 230, 229, 229, 228, 230, 230, 231, 230, 229, 230, 231, 231, 230, 229, 230, 230, 231, 230, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 232, 231, 230, 230, 232, 231, 231, 231, 230, 230, 232, 231, 230, 230, 230, 231, 231, 232, 231, 230, 231, 231, 231, 231, 231, 230, 231, 231, 231, 231, 230, 231, 232, 231, 231, 231, 231, 232, 232, 232, 231, 232, 232, 233, 233, 232, 232, 232, 234, 233, 234, 234, 233, 233, 232, 218, 188, 184, 188, 190, 184, 189, 188, 181, 177, 178, 179, 183, 185, 188, 186, 188, 183, 188, 191, 201, 212, 224, 222, 193, 217, 205, 102, 39, 36, 39, 47, 100, 130, 94, 88, 101, 69, 40, 41, 39, 39, 39, 44, 41, 43, 44, 37, 40, 52, 47, 49, 50, 68, 60, 61, 144, 156, 80, 49, 47, 54, 47, 51, 50, 45, 49, 53, 55, 77, 131, 159, 103, 55, 52, 67, 73, 88, 139, 229, 234, 233, 227, 206, 148, 93, 67, 75, 98, 131, 172, 224, 230, 231, 230, 230, 229, 228, 230, 230, 231, 230, 230, 230, 231, 231, 231, 229, 231, 230, 230, 230, 229, 228, 228, 230, 230, 229, 228, 229, 227, 222, 226, 221, 217, 223, 123, 220, 228, 227, 227, 224, 227, 228, 228, 228, 226, 225, 225, 227, 228, 227, 228, 228, 229, 230, 229, 229, 228, 229, 229, 230, 228, 228, 229, 230, 231, 230, 229, 229, 229, 230, 231, 229, 229, 229, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 229, 229, 231, 232, 231, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 231, 230, 230, 231, 231, 232, 230, 230, 230, 232, 232, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 231, 230, 230, 231, 232, 232, 231, 231, 230, 232, 232, 232, 231, 231, 232, 233, 233, 232, 233, 232, 234, 234, 233, 233, 233, 233, 232, 221, 197, 181, 188, 190, 183, 191, 191, 181, 180, 176, 181, 184, 187, 188, 185, 186, 183, 186, 186, 199, 207, 221, 224, 202, 204, 220, 145, 41, 38, 48, 60, 153, 80, 48, 49, 73, 134, 45, 41, 37, 38, 39, 39, 42, 40, 44, 43, 40, 61, 53, 42, 46, 46, 57, 63, 96, 157, 129, 53, 46, 51, 47, 47, 48, 48, 51, 56, 56, 102, 119, 162, 99, 57, 52, 63, 69, 94, 157, 231, 233, 232, 228, 199, 145, 83, 70, 83, 107, 138, 181, 225, 230, 231, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 229, 230, 230, 229, 229, 228, 229, 230, 231, 230, 228, 228, 227, 222, 224, 221, 220, 223, 124, 220, 227, 226, 226, 226, 228, 228, 228, 227, 226, 226, 227, 228, 227, 227, 228, 229, 229, 229, 230, 229, 229, 230, 230, 232, 229, 227, 229, 230, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 231, 230, 230, 230, 230, 230, 232, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 232, 231, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 232, 230, 230, 229, 231, 231, 231, 230, 230, 230, 232, 232, 231, 231, 230, 232, 232, 232, 231, 232, 232, 233, 233, 232, 232, 233, 234, 234, 234, 233, 234, 233, 232, 223, 201, 185, 184, 190, 184, 190, 189, 186, 185, 177, 178, 184, 188, 189, 183, 184, 176, 173, 181, 196, 206, 216, 225, 211, 188, 223, 170, 63, 45, 52, 72, 161, 105, 47, 52, 61, 148, 46, 37, 37, 38, 36, 37, 43, 44, 40, 42, 36, 43, 40, 42, 41, 56, 74, 63, 61, 141, 155, 71, 48, 49, 56, 50, 46, 51, 50, 63, 75, 106, 105, 164, 114, 62, 54, 70, 74, 97, 176, 232, 233, 232, 227, 199, 150, 84, 76, 87, 118, 135, 187, 226, 230, 231, 231, 231, 230, 230, 230, 231, 231, 229, 230, 230, 230, 231, 231, 230, 230, 230, 230, 229, 229, 228, 230, 230, 231, 231, 229, 229, 227, 222, 226, 221, 221, 223, 126, 219, 225, 227, 224, 227, 225, 229, 227, 226, 228, 227, 228, 229, 228, 228, 229, 229, 229, 229, 230, 229, 230, 230, 230, 230, 229, 229, 230, 230, 230, 230, 229, 229, 230, 230, 231, 230, 230, 229, 231, 231, 231, 230, 230, 230, 231, 230, 230, 229, 229, 231, 231, 231, 229, 229, 230, 231, 231, 231, 229, 230, 231, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 230, 229, 231, 231, 231, 231, 230, 230, 230, 232, 231, 231, 230, 230, 232, 232, 231, 230, 229, 230, 232, 232, 230, 230, 229, 231, 232, 231, 230, 230, 231, 231, 232, 231, 231, 231, 232, 232, 232, 231, 231, 232, 233, 233, 232, 233, 232, 233, 234, 234, 233, 234, 233, 233, 227, 200, 187, 184, 189, 186, 188, 190, 186, 179, 177, 178, 176, 179, 179, 178, 172, 173, 168, 174, 189, 204, 216, 228, 217, 187, 207, 195, 101, 41, 46, 61, 162, 166, 120, 78, 111, 109, 39, 37, 42, 37, 32, 37, 34, 41, 41, 43, 49, 79, 84, 48, 44, 69, 87, 66, 72, 119, 161, 125, 67, 52, 48, 48, 48, 51, 56, 61, 117, 87, 88, 169, 127, 58, 57, 66, 76, 99, 196, 232, 232, 231, 226, 195, 151, 83, 78, 102, 119, 144, 198, 227, 230, 231, 231, 231, 230, 229, 231, 231, 232, 229, 230, 231, 231, 231, 230, 230, 230, 230, 230, 230, 229, 229, 229, 229, 230, 230, 229, 228, 227, 222, 226, 220, 221, 224, 125, 217, 225, 227, 225, 227, 226, 229, 227, 228, 227, 227, 229, 228, 228, 228, 228, 229, 229, 229, 229, 228, 228, 230, 231, 231, 230, 229, 229, 230, 229, 231, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 230, 230, 230, 229, 229, 230, 231, 231, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 232, 230, 230, 230, 231, 231, 231, 230, 229, 231, 231, 231, 230, 230, 230, 231, 232, 232, 231, 230, 231, 231, 232, 230, 229, 230, 231, 231, 231, 231, 230, 231, 232, 232, 231, 230, 231, 232, 232, 232, 231, 231, 232, 233, 233, 232, 233, 233, 233, 234, 235, 234, 234, 234, 232, 230, 198, 180, 180, 188, 188, 186, 192, 188, 181, 169, 172, 174, 169, 174, 172, 169, 170, 169, 173, 181, 200, 214, 224, 225, 195, 194, 205, 143, 47, 41, 50, 104, 171, 173, 164, 136, 67, 43, 39, 39, 36, 38, 46, 40, 40, 37, 39, 38, 51, 50, 40, 44, 53, 61, 52, 61, 73, 164, 163, 138, 55, 49, 42, 46, 52, 56, 75, 145, 83, 76, 161, 139, 59, 56, 64, 81, 101, 214, 233, 232, 230, 225, 185, 142, 77, 80, 113, 132, 149, 209, 228, 230, 231, 231, 230, 230, 229, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 229, 230, 229, 228, 228, 228, 230, 231, 231, 229, 229, 227, 222, 229, 221, 222, 224, 120, 216, 226, 227, 225, 227, 228, 229, 229, 227, 227, 227, 229, 227, 229, 229, 228, 228, 229, 229, 230, 228, 227, 230, 230, 230, 230, 228, 229, 231, 230, 230, 229, 229, 229, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 228, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 231, 230, 230, 230, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 232, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 232, 231, 231, 230, 232, 232, 232, 231, 232, 231, 232, 233, 232, 232, 232, 234, 234, 235, 234, 234, 234, 233, 231, 197, 185, 181, 189, 191, 188, 191, 190, 181, 171, 169, 164, 166, 166, 170, 171, 175, 170, 172, 177, 193, 209, 219, 222, 207, 183, 203, 177, 85, 44, 53, 136, 119, 124, 168, 172, 156, 92, 43, 34, 36, 33, 62, 43, 40, 42, 44, 42, 36, 43, 38, 41, 45, 40, 47, 56, 81, 164, 169, 133, 49, 45, 44, 51, 55, 61, 122, 159, 78, 72, 157, 143, 66, 80, 68, 92, 122, 225, 233, 231, 228, 221, 174, 129, 81, 97, 114, 133, 151, 211, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 231, 230, 231, 231, 231, 230, 229, 229, 230, 229, 228, 229, 227, 231, 231, 229, 229, 230, 228, 221, 226, 224, 223, 224, 127, 220, 225, 226, 225, 228, 227, 228, 229, 228, 226, 227, 228, 228, 229, 227, 228, 228, 229, 230, 229, 228, 228, 228, 230, 230, 229, 228, 229, 230, 230, 231, 229, 229, 229, 231, 231, 230, 230, 230, 231, 231, 231, 229, 229, 230, 231, 231, 230, 230, 229, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 232, 232, 231, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 231, 230, 231, 231, 232, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 230, 228, 230, 231, 231, 231, 231, 230, 230, 232, 232, 231, 231, 231, 232, 232, 232, 231, 232, 232, 232, 233, 233, 232, 232, 233, 234, 234, 234, 234, 234, 234, 232, 211, 188, 181, 186, 192, 190, 195, 191, 190, 181, 167, 162, 160, 170, 166, 168, 173, 170, 166, 177, 189, 206, 212, 221, 216, 193, 192, 200, 139, 54, 100, 151, 52, 54, 70, 118, 159, 151, 49, 38, 40, 39, 40, 38, 36, 39, 42, 45, 38, 74, 38, 46, 39, 42, 47, 53, 87, 124, 185, 181, 60, 53, 53, 55, 58, 67, 139, 143, 86, 76, 154, 154, 94, 85, 76, 92, 162, 229, 232, 231, 227, 213, 166, 119, 85, 105, 120, 136, 156, 218, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 231, 229, 231, 231, 230, 230, 229, 229, 230, 229, 227, 229, 228, 231, 231, 230, 230, 230, 227, 222, 229, 226, 221, 223, 121, 216, 225, 226, 226, 227, 228, 229, 229, 228, 228, 227, 229, 229, 227, 228, 228, 228, 229, 230, 229, 228, 229, 228, 230, 230, 229, 229, 229, 230, 231, 231, 229, 230, 230, 231, 231, 230, 230, 229, 230, 230, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 231, 229, 229, 230, 231, 231, 231, 230, 230, 230, 231, 232, 231, 231, 231, 232, 232, 232, 232, 231, 232, 233, 233, 232, 232, 232, 233, 234, 234, 234, 234, 234, 234, 232, 222, 196, 183, 186, 188, 189, 193, 193, 194, 183, 169, 162, 163, 168, 171, 167, 169, 166, 172, 175, 179, 199, 211, 215, 219, 206, 185, 212, 178, 90, 115, 148, 43, 43, 41, 53, 104, 162, 66, 41, 42, 45, 46, 46, 46, 42, 41, 39, 38, 41, 47, 48, 44, 60, 40, 57, 52, 59, 163, 205, 113, 71, 68, 76, 79, 82, 81, 63, 58, 56, 148, 156, 68, 65, 78, 105, 190, 232, 231, 230, 226, 195, 159, 98, 103, 115, 124, 138, 176, 221, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 230, 231, 231, 229, 229, 229, 230, 230, 229, 228, 229, 230, 231, 229, 229, 230, 227, 222, 228, 222, 218, 224, 117, 220, 226, 226, 227, 225, 227, 229, 228, 227, 227, 226, 228, 228, 228, 227, 227, 228, 229, 230, 229, 229, 228, 229, 230, 230, 229, 229, 229, 230, 230, 230, 230, 229, 230, 231, 231, 229, 229, 230, 231, 230, 230, 229, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 229, 229, 230, 231, 232, 231, 230, 230, 231, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 230, 230, 230, 231, 231, 230, 229, 230, 230, 231, 232, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 232, 231, 231, 230, 232, 232, 232, 231, 231, 232, 233, 233, 233, 232, 232, 233, 234, 234, 233, 234, 234, 234, 232, 227, 206, 185, 180, 190, 192, 194, 197, 196, 185, 171, 164, 161, 164, 175, 168, 172, 162, 164, 169, 172, 189, 202, 208, 218, 213, 193, 197, 195, 144, 95, 149, 56, 34, 38, 48, 70, 155, 58, 80, 137, 142, 149, 142, 138, 135, 104, 35, 35, 39, 52, 61, 34, 66, 42, 67, 43, 61, 96, 204, 173, 149, 167, 163, 168, 160, 143, 56, 53, 55, 140, 164, 69, 64, 110, 184, 223, 232, 231, 227, 224, 182, 147, 94, 110, 123, 134, 146, 190, 224, 230, 230, 231, 230, 230, 230, 229, 231, 231, 231, 230, 230, 230, 231, 231, 231, 229, 229, 229, 230, 231, 228, 228, 229, 230, 231, 230, 230, 230, 227, 222, 228, 222, 222, 224, 119, 217, 225, 226, 227, 226, 227, 228, 228, 227, 228, 227, 228, 229, 230, 228, 227, 227, 229, 229, 230, 228, 228, 229, 230, 231, 229, 229, 229, 230, 231, 231, 230, 230, 229, 231, 230, 230, 229, 230, 231, 230, 230, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 229, 229, 230, 231, 232, 230, 230, 230, 231, 232, 231, 230, 230, 230, 232, 231, 231, 230, 230, 231, 231, 231, 231, 230, 230, 231, 231, 231, 229, 230, 230, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 230, 232, 232, 232, 231, 231, 232, 233, 232, 232, 232, 232, 233, 234, 234, 233, 234, 234, 235, 233, 230, 211, 185, 177, 188, 193, 192, 195, 200, 191, 177, 164, 162, 170, 174, 177, 169, 169, 157, 145, 173, 177, 191, 205, 221, 218, 202, 182, 196, 177, 98, 125, 114, 50, 38, 44, 103, 105, 46, 122, 173, 179, 182, 180, 174, 164, 92, 40, 42, 41, 42, 39, 43, 63, 51, 46, 39, 51, 62, 169, 201, 152, 156, 149, 150, 133, 105, 50, 51, 58, 120, 137, 66, 71, 95, 172, 229, 232, 231, 226, 214, 173, 131, 98, 116, 124, 135, 144, 205, 227, 230, 230, 231, 231, 230, 230, 230, 230, 231, 232, 230, 230, 230, 231, 231, 230, 228, 228, 228, 230, 231, 229, 229, 228, 230, 231, 231, 229, 229, 228, 223, 228, 224, 222, 226, 114, 217, 225, 226, 228, 226, 228, 226, 227, 227, 227, 228, 228, 229, 230, 228, 227, 227, 230, 230, 230, 228, 228, 229, 230, 229, 229, 228, 229, 231, 230, 231, 229, 230, 230, 231, 231, 230, 229, 229, 231, 231, 230, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 230, 231, 230, 230, 229, 229, 231, 231, 231, 230, 230, 232, 232, 231, 230, 230, 231, 231, 231, 231, 230, 230, 231, 231, 231, 231, 230, 231, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 231, 231, 229, 232, 232, 232, 231, 231, 231, 232, 232, 232, 232, 232, 232, 234, 234, 233, 233, 234, 234, 234, 230, 214, 185, 184, 188, 191, 191, 200, 205, 191, 182, 167, 166, 166, 177, 186, 175, 174, 173, 164, 176, 181, 186, 202, 213, 218, 210, 190, 187, 186, 145, 70, 94, 89, 70, 71, 72, 43, 43, 84, 93, 100, 100, 98, 98, 142, 48, 41, 41, 38, 46, 89, 119, 98, 127, 118, 59, 50, 59, 119, 198, 135, 70, 79, 73, 62, 53, 49, 43, 48, 52, 58, 63, 73, 94, 204, 231, 230, 228, 222, 198, 159, 114, 107, 120, 130, 136, 162, 216, 229, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 231, 230, 230, 231, 231, 230, 229, 229, 228, 230, 230, 228, 229, 229, 231, 231, 231, 230, 229, 227, 222, 226, 223, 222, 224, 116, 214, 225, 226, 226, 225, 224, 228, 228, 228, 226, 227, 228, 230, 230, 229, 228, 229, 229, 230, 230, 227, 228, 229, 230, 230, 229, 228, 230, 231, 230, 231, 229, 230, 229, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 229, 229, 230, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 231, 230, 231, 230, 230, 230, 231, 231, 231, 231, 230, 230, 232, 232, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 231, 230, 230, 230, 230, 232, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 230, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 232, 232, 233, 234, 234, 233, 233, 233, 235, 233, 230, 222, 181, 182, 181, 192, 194, 194, 201, 194, 185, 171, 167, 167, 178, 187, 184, 181, 178, 181, 183, 189, 183, 193, 206, 215, 216, 208, 181, 196, 175, 114, 47, 41, 41, 36, 36, 38, 35, 38, 37, 38, 46, 53, 119, 112, 39, 37, 44, 48, 91, 140, 60, 52, 75, 145, 131, 51, 50, 64, 163, 149, 104, 95, 107, 127, 83, 54, 42, 49, 50, 54, 65, 83, 146, 222, 232, 230, 224, 217, 173, 141, 118, 116, 126, 128, 139, 182, 224, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 230, 230, 230, 230, 230, 230, 230, 229, 229, 230, 230, 228, 229, 229, 231, 231, 230, 228, 229, 227, 223, 227, 225, 222, 224, 113, 210, 227, 226, 225, 222, 226, 228, 228, 226, 228, 227, 227, 229, 229, 228, 227, 228, 229, 229, 230, 228, 228, 229, 229, 230, 228, 228, 230, 231, 230, 230, 230, 229, 230, 231, 230, 229, 230, 229, 231, 231, 230, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 231, 230, 230, 230, 231, 232, 231, 229, 230, 230, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 232, 231, 231, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 233, 233, 233, 233, 233, 233, 234, 234, 232, 228, 186, 181, 185, 186, 195, 192, 197, 199, 192, 176, 166, 162, 177, 188, 185, 184, 185, 186, 183, 191, 187, 188, 199, 211, 212, 215, 189, 185, 194, 159, 79, 42, 37, 37, 33, 36, 34, 38, 38, 43, 52, 81, 156, 74, 35, 36, 53, 58, 147, 121, 43, 48, 47, 106, 114, 48, 46, 47, 58, 95, 50, 51, 58, 108, 151, 84, 45, 51, 48, 58, 75, 88, 197, 228, 230, 228, 224, 194, 157, 127, 117, 117, 122, 129, 147, 201, 228, 229, 230, 230, 231, 232, 231, 230, 230, 231, 232, 231, 229, 230, 229, 230, 230, 230, 230, 230, 229, 229, 228, 229, 229, 229, 230, 230, 230, 230, 229, 227, 224, 225, 225, 223, 223, 114, 213, 226, 227, 224, 224, 225, 227, 227, 226, 227, 228, 228, 229, 228, 227, 228, 228, 230, 230, 230, 229, 230, 229, 229, 230, 230, 229, 229, 230, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 230, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 229, 231, 231, 231, 230, 230, 230, 231, 231, 231, 229, 230, 231, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 232, 230, 230, 231, 232, 233, 231, 231, 231, 232, 233, 233, 233, 232, 234, 234, 234, 232, 227, 204, 178, 183, 189, 193, 190, 192, 196, 193, 183, 170, 170, 178, 186, 183, 183, 184, 190, 185, 184, 190, 180, 189, 206, 204, 205, 206, 184, 188, 184, 146, 63, 38, 37, 32, 35, 38, 35, 35, 40, 55, 134, 156, 48, 37, 40, 50, 89, 168, 93, 40, 41, 45, 52, 48, 41, 42, 40, 53, 97, 43, 45, 56, 67, 155, 137, 51, 48, 56, 60, 82, 140, 223, 227, 228, 225, 217, 170, 142, 121, 121, 118, 124, 137, 168, 217, 230, 230, 229, 230, 232, 231, 231, 230, 230, 230, 231, 231, 229, 229, 230, 231, 230, 230, 229, 229, 227, 229, 229, 228, 227, 228, 230, 229, 230, 228, 229, 226, 222, 229, 225, 222, 224, 121, 214, 226, 227, 227, 226, 227, 228, 227, 228, 228, 227, 228, 230, 228, 227, 228, 227, 230, 229, 230, 230, 229, 228, 229, 230, 230, 229, 229, 230, 230, 231, 230, 229, 230, 231, 231, 230, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 231, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 229, 230, 231, 230, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 231, 230, 230, 229, 231, 231, 230, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 231, 231, 230, 231, 231, 232, 231, 231, 230, 231, 232, 233, 232, 232, 231, 233, 234, 233, 233, 233, 233, 235, 235, 233, 228, 223, 177, 185, 183, 194, 191, 193, 199, 193, 189, 176, 168, 174, 181, 182, 186, 189, 190, 192, 191, 189, 189, 182, 191, 202, 206, 211, 197, 176, 192, 176, 131, 50, 39, 35, 36, 35, 36, 39, 51, 68, 165, 137, 37, 35, 39, 47, 123, 166, 77, 42, 61, 84, 98, 63, 41, 41, 47, 104, 115, 40, 42, 51, 57, 145, 158, 67, 52, 62, 71, 101, 203, 227, 226, 227, 224, 192, 161, 127, 122, 118, 118, 123, 137, 191, 226, 231, 229, 229, 229, 230, 231, 230, 230, 230, 230, 232, 230, 230, 229, 228, 230, 230, 230, 229, 228, 227, 229, 228, 228, 228, 227, 228, 229, 229, 229, 229, 225, 221, 227, 224, 223, 225, 131, 213, 225, 229, 225, 225, 226, 227, 228, 228, 228, 227, 227, 229, 228, 227, 226, 225, 225, 228, 228, 228, 229, 228, 229, 229, 229, 229, 228, 230, 230, 230, 230, 229, 230, 231, 231, 230, 228, 229, 230, 231, 231, 229, 229, 229, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 229, 229, 230, 231, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 229, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 231, 232, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 232, 231, 233, 233, 233, 232, 232, 233, 234, 235, 233, 231, 228, 191, 180, 186, 184, 192, 192, 192, 192, 193, 179, 173, 175, 182, 184, 184, 189, 186, 189, 186, 189, 188, 184, 182, 196, 208, 211, 208, 191, 178, 189, 172, 114, 47, 37, 37, 34, 41, 35, 47, 108, 165, 109, 37, 34, 38, 46, 132, 165, 72, 54, 67, 73, 121, 142, 102, 43, 45, 115, 84, 40, 41, 49, 55, 143, 160, 69, 54, 64, 86, 173, 221, 226, 225, 225, 210, 175, 133, 121, 119, 115, 117, 123, 158, 209, 229, 230, 230, 229, 228, 230, 231, 230, 229, 230, 229, 232, 231, 229, 229, 227, 229, 230, 230, 229, 228, 228, 228, 229, 227, 225, 225, 228, 228, 227, 229, 228, 224, 220, 227, 224, 224, 224, 126, 214, 226, 228, 225, 227, 227, 227, 229, 229, 228, 227, 227, 229, 228, 226, 223, 224, 227, 228, 228, 228, 227, 227, 227, 228, 228, 227, 229, 230, 230, 229, 230, 229, 230, 230, 230, 230, 230, 230, 230, 231, 231, 229, 229, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 231, 232, 231, 231, 230, 230, 230, 231, 231, 230, 231, 231, 231, 231, 231, 231, 231, 231, 232, 232, 231, 231, 231, 232, 233, 232, 231, 231, 232, 233, 233, 233, 233, 232, 234, 234, 234, 232, 228, 217, 177, 185, 182, 191, 191, 192, 198, 192, 188, 175, 173, 179, 182, 184, 186, 188, 184, 187, 187, 184, 186, 178, 186, 202, 205, 209, 203, 183, 179, 193, 163, 109, 42, 35, 35, 39, 41, 43, 141, 169, 96, 34, 37, 40, 49, 136, 166, 84, 56, 42, 44, 53, 135, 158, 77, 50, 92, 94, 41, 41, 50, 54, 142, 160, 69, 62, 76, 138, 216, 227, 225, 224, 218, 177, 158, 121, 111, 112, 106, 107, 126, 180, 220, 230, 231, 229, 228, 229, 230, 231, 230, 229, 229, 229, 230, 231, 228, 229, 227, 228, 229, 228, 228, 226, 225, 228, 228, 226, 224, 225, 227, 229, 229, 228, 227, 224, 219, 225, 225, 224, 225, 135, 220, 227, 225, 225, 227, 228, 228, 229, 230, 229, 227, 226, 228, 227, 224, 223, 224, 224, 228, 229, 227, 224, 226, 225, 224, 225, 227, 228, 230, 230, 228, 229, 229, 230, 230, 230, 230, 230, 230, 231, 231, 231, 229, 229, 229, 231, 231, 231, 229, 230, 231, 232, 231, 230, 230, 230, 231, 231, 231, 229, 230, 230, 230, 231, 230, 230, 230, 230, 231, 232, 230, 230, 230, 231, 230, 229, 229, 230, 230, 230, 230, 230, 230, 230, 232, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 231, 230, 230, 232, 232, 231, 230, 230, 232, 232, 231, 230, 231, 231, 232, 232, 232, 231, 231, 233, 233, 233, 233, 232, 233, 234, 234, 234, 231, 230, 227, 187, 183, 183, 187, 187, 195, 189, 192, 190, 182, 171, 178, 178, 180, 187, 187, 185, 187, 192, 185, 185, 181, 173, 193, 204, 209, 208, 201, 179, 184, 189, 162, 100, 42, 36, 36, 44, 46, 154, 167, 73, 37, 33, 41, 48, 132, 169, 87, 59, 36, 41, 46, 94, 161, 123, 45, 50, 98, 41, 41, 56, 71, 154, 129, 58, 73, 119, 208, 224, 226, 224, 220, 191, 165, 125, 111, 97, 103, 100, 109, 144, 211, 228, 231, 230, 229, 228, 229, 229, 229, 230, 228, 229, 228, 231, 229, 228, 227, 226, 229, 229, 227, 225, 224, 226, 226, 226, 225, 225, 226, 226, 226, 227, 226, 226, 222, 218, 227, 224, 222, 226, 127, 218, 228, 226, 225, 226, 227, 229, 229, 230, 228, 228, 227, 228, 225, 223, 221, 222, 223, 227, 227, 225, 224, 226, 226, 225, 225, 227, 226, 228, 227, 227, 227, 227, 229, 230, 231, 230, 229, 230, 231, 231, 231, 229, 229, 229, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 230, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 230, 229, 230, 230, 230, 231, 229, 229, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 231, 229, 230, 231, 231, 231, 230, 230, 230, 231, 232, 231, 231, 230, 231, 231, 231, 231, 231, 231, 232, 232, 232, 231, 232, 233, 233, 233, 232, 232, 233, 234, 234, 233, 232, 231, 228, 212, 183, 184, 181, 186, 194, 191, 193, 194, 188, 174, 179, 180, 182, 184, 187, 186, 188, 186, 185, 178, 180, 168, 179, 194, 197, 207, 209, 199, 178, 174, 185, 159, 101, 47, 41, 48, 53, 159, 163, 68, 34, 37, 36, 50, 112, 160, 104, 60, 36, 37, 51, 72, 156, 144, 45, 41, 68, 90, 69, 70, 128, 135, 67, 71, 112, 196, 220, 223, 224, 219, 197, 164, 129, 116, 88, 87, 87, 89, 110, 179, 220, 229, 230, 230, 229, 228, 229, 229, 229, 230, 228, 228, 229, 230, 230, 227, 228, 228, 230, 225, 225, 222, 225, 227, 226, 227, 226, 224, 224, 227, 225, 225, 223, 222, 220, 215, 228, 224, 223, 223, 119, 217, 227, 227, 225, 227, 227, 229, 228, 229, 228, 226, 226, 227, 225, 220, 221, 224, 225, 225, 229, 226, 225, 226, 224, 226, 225, 225, 225, 227, 227, 228, 227, 229, 228, 228, 230, 230, 228, 228, 230, 230, 230, 229, 230, 230, 230, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 229, 230, 230, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 229, 230, 231, 230, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 232, 231, 230, 229, 231, 231, 232, 231, 230, 231, 232, 233, 231, 231, 231, 232, 233, 233, 232, 232, 233, 233, 233, 233, 232, 232, 230, 227, 180, 182, 177, 184, 194, 189, 197, 191, 189, 182, 176, 174, 178, 181, 183, 188, 186, 184, 181, 172, 165, 156, 163, 174, 192, 202, 203, 205, 193, 173, 182, 178, 163, 111, 54, 53, 58, 151, 150, 60, 34, 36, 37, 52, 86, 157, 118, 74, 40, 40, 48, 60, 160, 149, 42, 38, 40, 50, 72, 77, 82, 84, 151, 117, 194, 218, 218, 220, 216, 196, 171, 128, 112, 90, 79, 76, 82, 91, 145, 206, 225, 230, 230, 230, 229, 228, 229, 230, 229, 229, 227, 229, 230, 230, 230, 226, 228, 227, 229, 225, 227, 226, 226, 225, 225, 226, 226, 223, 223, 226, 223, 225, 224, 222, 220, 214, 226, 224, 221, 225, 118, 220, 227, 227, 226, 229, 227, 227, 229, 228, 228, 226, 227, 224, 222, 217, 218, 220, 224, 225, 228, 225, 226, 224, 225, 224, 224, 226, 227, 226, 227, 228, 226, 229, 227, 228, 229, 229, 228, 229, 230, 228, 229, 229, 229, 229, 230, 230, 231, 229, 229, 230, 230, 231, 230, 230, 229, 231, 231, 229, 229, 229, 230, 230, 231, 229, 229, 230, 231, 231, 230, 230, 229, 230, 230, 230, 229, 229, 229, 230, 229, 229, 228, 228, 229, 230, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 232, 231, 230, 230, 231, 231, 231, 231, 230, 231, 232, 232, 232, 231, 231, 233, 233, 232, 232, 232, 232, 232, 233, 233, 233, 233, 232, 230, 205, 177, 182, 178, 191, 195, 193, 187, 190, 188, 181, 168, 175, 178, 179, 187, 187, 185, 176, 162, 154, 151, 154, 162, 178, 190, 202, 208, 203, 192, 171, 175, 183, 166, 134, 111, 82, 57, 53, 40, 32, 34, 36, 51, 53, 142, 142, 74, 56, 44, 49, 57, 155, 129, 37, 40, 39, 36, 43, 46, 58, 102, 188, 200, 213, 219, 215, 216, 194, 173, 142, 104, 99, 69, 73, 74, 80, 117, 188, 221, 228, 230, 230, 230, 229, 229, 229, 230, 228, 229, 228, 229, 229, 230, 229, 227, 227, 226, 228, 224, 227, 225, 227, 226, 227, 227, 226, 222, 222, 225, 224, 226, 224, 223, 221, 214, 226, 224, 221, 224, 121, 219, 225, 225, 227, 227, 227, 229, 230, 226, 226, 224, 226, 224, 226, 218, 217, 220, 224, 224, 225, 224, 224, 225, 226, 225, 223, 227, 225, 227, 228, 227, 227, 227, 227, 228, 229, 229, 229, 229, 230, 229, 230, 228, 229, 229, 229, 231, 230, 229, 229, 230, 230, 229, 229, 229, 228, 229, 228, 227, 226, 227, 227, 227, 227, 224, 226, 224, 224, 223, 220, 218, 217, 214, 217, 210, 206, 208, 203, 198, 199, 196, 189, 189, 190, 199, 219, 221, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 231, 230, 231, 231, 231, 231, 230, 230, 231, 231, 231, 231, 231, 231, 232, 232, 231, 231, 231, 232, 233, 233, 232, 232, 232, 233, 234, 234, 233, 233, 232, 230, 227, 171, 176, 179, 184, 193, 193, 186, 188, 186, 185, 175, 167, 174, 178, 185, 184, 179, 176, 153, 149, 149, 146, 146, 160, 175, 192, 199, 204, 199, 192, 168, 176, 183, 177, 153, 103, 50, 43, 41, 35, 36, 38, 44, 52, 99, 137, 85, 57, 41, 52, 72, 153, 77, 34, 38, 35, 36, 44, 54, 78, 157, 205, 215, 215, 210, 205, 189, 164, 129, 105, 91, 74, 68, 65, 74, 96, 166, 215, 227, 229, 231, 230, 230, 228, 228, 229, 229, 229, 229, 228, 229, 229, 230, 227, 228, 227, 226, 226, 227, 227, 224, 227, 228, 229, 228, 226, 225, 224, 224, 225, 224, 225, 223, 220, 212, 229, 226, 223, 227, 131, 223, 225, 228, 227, 228, 229, 231, 231, 228, 223, 210, 203, 198, 202, 193, 194, 193, 195, 196, 196, 194, 196, 193, 196, 197, 197, 200, 197, 200, 204, 199, 202, 206, 204, 206, 206, 208, 210, 211, 211, 212, 219, 214, 215, 218, 218, 226, 212, 203, 201, 198, 193, 189, 186, 182, 178, 169, 166, 159, 160, 163, 157, 152, 156, 148, 148, 136, 138, 134, 133, 133, 128, 122, 126, 116, 117, 116, 111, 111, 115, 120, 124, 124, 132, 154, 132, 140, 226, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 231, 231, 230, 230, 231, 232, 231, 231, 231, 231, 232, 232, 231, 231, 231, 232, 233, 232, 231, 232, 232, 233, 234, 234, 233, 234, 234, 233, 228, 201, 172, 178, 182, 190, 189, 185, 185, 188, 184, 181, 173, 164, 175, 182, 183, 184, 171, 153, 146, 142, 135, 139, 140, 150, 171, 189, 193, 199, 203, 190, 172, 172, 186, 186, 167, 123, 68, 50, 42, 39, 44, 39, 46, 66, 98, 131, 62, 48, 51, 109, 118, 39, 37, 36, 39, 43, 59, 111, 175, 202, 208, 209, 206, 199, 178, 161, 130, 105, 100, 66, 69, 71, 62, 85, 143, 203, 226, 228, 229, 230, 231, 229, 229, 229, 230, 230, 230, 228, 229, 228, 227, 228, 228, 228, 227, 227, 227, 225, 223, 224, 226, 226, 227, 228, 224, 226, 225, 225, 224, 225, 225, 221, 218, 214, 233, 229, 226, 231, 134, 226, 234, 235, 235, 237, 237, 240, 238, 227, 204, 95, 91, 82, 80, 81, 81, 80, 85, 85, 85, 79, 82, 80, 81, 78, 82, 79, 77, 81, 83, 84, 81, 81, 82, 87, 86, 81, 88, 87, 92, 94, 103, 97, 101, 108, 127, 160, 143, 124, 131, 133, 124, 110, 109, 104, 97, 96, 99, 96, 95, 95, 92, 95, 99, 97, 93, 88, 95, 96, 93, 91, 90, 94, 89, 91, 91, 94, 97, 103, 107, 111, 112, 114, 110, 151, 106, 117, 225, 230, 231, 230, 231, 229, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 230, 232, 232, 230, 230, 231, 232, 232, 232, 231, 231, 232, 233, 232, 232, 232, 232, 234, 234, 233, 233, 233, 235, 233, 230, 224, 171, 178, 183, 182, 187, 191, 186, 188, 189, 187, 180, 168, 162, 167, 173, 173, 161, 139, 140, 131, 127, 131, 127, 138, 143, 171, 182, 188, 200, 199, 195, 177, 161, 176, 187, 177, 159, 108, 58, 45, 38, 48, 46, 52, 55, 95, 111, 96, 82, 93, 54, 55, 77, 90, 65, 97, 154, 187, 201, 201, 201, 201, 182, 170, 155, 125, 107, 100, 64, 59, 67, 69, 76, 131, 193, 221, 229, 229, 230, 231, 231, 230, 230, 229, 229, 230, 231, 230, 230, 228, 228, 230, 228, 225, 228, 227, 226, 225, 225, 223, 225, 227, 228, 225, 225, 226, 225, 224, 226, 223, 223, 223, 218, 215, 235, 229, 228, 232, 123, 226, 233, 232, 235, 236, 238, 240, 238, 228, 203, 84, 80, 70, 75, 72, 71, 69, 73, 76, 75, 71, 74, 72, 74, 72, 66, 67, 70, 69, 72, 75, 71, 76, 73, 75, 74, 73, 74, 70, 76, 78, 79, 75, 80, 99, 139, 158, 159, 130, 143, 121, 109, 95, 87, 92, 86, 86, 89, 88, 95, 86, 86, 90, 92, 89, 90, 86, 88, 91, 90, 79, 83, 80, 87, 86, 90, 95, 104, 112, 116, 124, 120, 146, 106, 145, 105, 118, 224, 230, 231, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 232, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 232, 232, 232, 233, 234, 233, 233, 233, 235, 235, 234, 229, 204, 177, 178, 187, 187, 190, 189, 187, 188, 188, 190, 178, 170, 155, 153, 148, 142, 143, 137, 132, 140, 123, 122, 121, 128, 138, 162, 174, 184, 191, 200, 195, 183, 163, 162, 178, 182, 171, 150, 110, 79, 95, 93, 88, 88, 84, 71, 170, 97, 109, 113, 131, 132, 138, 151, 175, 188, 190, 197, 191, 182, 174, 167, 146, 108, 120, 97, 64, 53, 61, 62, 75, 121, 185, 222, 230, 230, 229, 230, 231, 231, 230, 229, 229, 230, 231, 230, 229, 229, 228, 230, 229, 230, 226, 227, 228, 224, 225, 224, 224, 224, 228, 226, 226, 226, 225, 226, 226, 224, 222, 223, 221, 219, 213, 234, 229, 230, 230, 127, 224, 230, 233, 234, 235, 237, 241, 238, 228, 202, 87, 79, 98, 74, 69, 70, 73, 72, 73, 77, 74, 74, 75, 74, 73, 70, 68, 72, 70, 71, 75, 73, 74, 80, 80, 83, 80, 83, 80, 84, 84, 82, 79, 84, 96, 148, 170, 179, 166, 207, 113, 115, 103, 89, 97, 113, 103, 102, 133, 160, 165, 165, 171, 174, 173, 154, 150, 153, 167, 131, 102, 140, 129, 131, 143, 153, 160, 169, 170, 178, 176, 160, 158, 105, 139, 101, 116, 222, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 231, 231, 231, 230, 232, 232, 231, 230, 230, 230, 232, 232, 232, 231, 231, 232, 232, 232, 231, 232, 232, 234, 234, 233, 233, 233, 235, 235, 234, 231, 227, 191, 174, 181, 183, 184, 191, 192, 187, 189, 189, 183, 173, 157, 147, 142, 136, 135, 135, 133, 132, 129, 123, 114, 113, 118, 134, 158, 167, 181, 192, 195, 199, 189, 169, 157, 160, 178, 180, 164, 159, 139, 119, 110, 105, 107, 108, 150, 117, 128, 139, 153, 161, 165, 169, 172, 174, 176, 175, 171, 165, 151, 126, 119, 118, 90, 62, 53, 56, 59, 73, 117, 180, 217, 229, 231, 230, 230, 229, 231, 230, 231, 229, 229, 230, 231, 230, 229, 229, 227, 227, 228, 228, 226, 227, 228, 226, 227, 226, 225, 224, 225, 224, 224, 225, 224, 223, 224, 225, 224, 223, 222, 219, 218, 231, 228, 227, 228, 120, 221, 229, 231, 231, 233, 235, 236, 232, 223, 190, 89, 78, 151, 75, 75, 82, 121, 130, 138, 144, 153, 156, 168, 164, 159, 142, 141, 148, 156, 146, 152, 153, 141, 186, 191, 192, 193, 195, 194, 197, 192, 181, 158, 95, 92, 136, 170, 190, 169, 212, 190, 211, 183, 153, 147, 177, 158, 146, 200, 223, 225, 225, 225, 222, 217, 184, 192, 171, 162, 127, 108, 150, 144, 148, 160, 170, 168, 177, 176, 183, 180, 163, 155, 104, 143, 102, 112, 223, 229, 232, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 228, 230, 231, 232, 231, 230, 230, 231, 232, 232, 232, 231, 231, 232, 233, 232, 232, 232, 232, 234, 234, 233, 233, 233, 234, 235, 235, 233, 230, 225, 177, 177, 179, 180, 187, 192, 190, 187, 192, 187, 185, 174, 159, 144, 137, 133, 135, 128, 129, 133, 120, 117, 89, 81, 110, 154, 147, 156, 175, 188, 198, 193, 190, 185, 166, 153, 154, 167, 172, 170, 168, 161, 154, 147, 142, 153, 147, 142, 152, 156, 156, 160, 165, 169, 174, 172, 170, 155, 129, 125, 131, 116, 80, 63, 69, 61, 56, 68, 124, 182, 217, 227, 230, 231, 230, 229, 229, 229, 229, 229, 229, 230, 229, 230, 229, 230, 228, 228, 227, 229, 228, 226, 228, 227, 225, 227, 226, 224, 227, 226, 226, 225, 227, 226, 225, 226, 223, 224, 224, 223, 221, 219, 231, 227, 227, 228, 122, 221, 231, 231, 230, 233, 233, 236, 232, 223, 190, 87, 88, 105, 85, 96, 103, 177, 181, 182, 186, 185, 185, 187, 185, 159, 137, 141, 139, 143, 142, 144, 158, 176, 219, 222, 223, 223, 220, 222, 223, 214, 201, 187, 107, 94, 150, 176, 178, 164, 201, 200, 222, 195, 182, 172, 192, 171, 160, 208, 229, 231, 231, 232, 227, 217, 172, 151, 100, 85, 78, 79, 95, 126, 146, 155, 168, 171, 177, 180, 183, 179, 156, 158, 104, 136, 97, 121, 225, 230, 231, 231, 231, 230, 230, 229, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 230, 230, 230, 231, 232, 232, 231, 230, 231, 232, 232, 231, 231, 231, 231, 231, 232, 232, 232, 232, 233, 233, 233, 232, 233, 234, 235, 235, 234, 233, 230, 223, 200, 183, 183, 181, 188, 194, 190, 188, 187, 184, 180, 170, 160, 151, 135, 132, 132, 126, 130, 125, 126, 113, 79, 161, 155, 109, 119, 144, 168, 181, 186, 189, 192, 194, 184, 165, 145, 140, 152, 166, 171, 169, 178, 169, 168, 168, 172, 172, 173, 176, 173, 172, 166, 161, 146, 131, 136, 135, 135, 109, 69, 83, 60, 54, 64, 77, 119, 184, 219, 227, 230, 230, 230, 229, 228, 228, 229, 231, 230, 229, 229, 229, 229, 230, 229, 229, 229, 230, 228, 228, 227, 226, 223, 224, 227, 228, 225, 226, 228, 225, 226, 225, 225, 225, 225, 223, 223, 220, 223, 220, 216, 232, 228, 227, 228, 132, 224, 230, 232, 231, 234, 235, 237, 233, 222, 187, 87, 74, 94, 112, 119, 121, 130, 129, 131, 136, 134, 135, 140, 143, 146, 148, 152, 152, 141, 115, 125, 140, 174, 220, 226, 224, 224, 222, 222, 223, 220, 204, 192, 110, 87, 124, 176, 157, 160, 183, 203, 223, 203, 185, 183, 195, 179, 173, 207, 231, 232, 233, 233, 227, 213, 143, 80, 78, 85, 85, 79, 85, 102, 145, 158, 166, 172, 174, 180, 181, 182, 156, 159, 116, 142, 102, 122, 226, 230, 231, 231, 231, 229, 230, 230, 231, 231, 230, 230, 229, 231, 231, 231, 230, 230, 231, 231, 232, 230, 230, 230, 232, 232, 232, 231, 230, 231, 232, 232, 231, 231, 231, 231, 232, 233, 231, 232, 232, 233, 233, 232, 232, 232, 234, 235, 235, 234, 234, 233, 232, 226, 189, 182, 184, 183, 192, 195, 188, 182, 188, 185, 179, 171, 157, 145, 137, 131, 131, 127, 121, 124, 119, 77, 167, 116, 71, 79, 110, 126, 153, 168, 178, 186, 189, 190, 188, 180, 174, 164, 152, 143, 135, 142, 151, 159, 159, 158, 156, 162, 155, 148, 139, 135, 142, 149, 147, 145, 118, 79, 54, 45, 64, 79, 57, 63, 81, 141, 212, 227, 230, 230, 231, 232, 230, 229, 229, 230, 231, 230, 230, 229, 230, 230, 229, 229, 229, 229, 230, 230, 228, 225, 225, 222, 226, 228, 228, 226, 227, 226, 226, 227, 226, 224, 224, 225, 224, 224, 223, 224, 220, 218, 232, 227, 228, 227, 133, 224, 232, 233, 232, 235, 236, 236, 233, 222, 178, 94, 74, 87, 117, 125, 122, 122, 126, 137, 134, 138, 139, 145, 150, 151, 148, 151, 133, 117, 107, 119, 132, 179, 221, 227, 225, 222, 224, 216, 220, 221, 194, 189, 104, 86, 116, 181, 145, 171, 186, 205, 228, 226, 213, 190, 201, 195, 183, 210, 232, 233, 235, 233, 228, 209, 119, 76, 77, 85, 81, 79, 82, 94, 119, 154, 172, 174, 172, 180, 185, 185, 161, 172, 114, 144, 101, 124, 226, 230, 231, 231, 230, 229, 229, 230, 231, 230, 230, 230, 230, 232, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 232, 231, 231, 231, 232, 232, 233, 231, 231, 231, 233, 233, 232, 232, 232, 234, 234, 235, 234, 234, 234, 235, 233, 226, 192, 180, 185, 185, 189, 193, 184, 182, 181, 187, 183, 172, 163, 149, 142, 139, 126, 124, 116, 99, 99, 105, 45, 56, 52, 86, 94, 100, 129, 147, 164, 175, 180, 180, 185, 188, 183, 189, 179, 176, 166, 162, 155, 151, 152, 151, 156, 161, 168, 161, 162, 161, 153, 130, 100, 71, 55, 42, 46, 69, 76, 75, 65, 70, 123, 202, 226, 229, 230, 231, 231, 229, 228, 229, 229, 231, 230, 230, 229, 229, 230, 230, 230, 229, 229, 229, 227, 225, 224, 223, 221, 225, 227, 227, 225, 226, 227, 226, 226, 226, 225, 224, 223, 224, 222, 222, 223, 219, 215, 231, 228, 227, 228, 116, 218, 232, 232, 233, 234, 236, 236, 234, 222, 178, 89, 78, 81, 116, 127, 128, 128, 140, 141, 135, 138, 138, 147, 150, 144, 123, 91, 78, 83, 87, 100, 130, 184, 223, 224, 224, 224, 220, 220, 222, 216, 208, 194, 99, 92, 124, 200, 147, 171, 181, 214, 230, 230, 227, 220, 211, 205, 195, 219, 232, 233, 235, 233, 224, 207, 115, 91, 92, 87, 81, 74, 79, 83, 99, 151, 166, 178, 179, 182, 189, 184, 158, 173, 123, 150, 107, 122, 225, 230, 231, 231, 230, 229, 229, 230, 230, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 231, 231, 231, 231, 232, 232, 233, 232, 231, 231, 232, 233, 233, 232, 232, 233, 234, 234, 233, 234, 234, 235, 235, 233, 228, 203, 184, 191, 185, 182, 186, 182, 176, 182, 179, 181, 174, 164, 154, 140, 127, 120, 116, 96, 172, 71, 52, 94, 104, 102, 95, 88, 90, 98, 116, 135, 150, 163, 168, 175, 180, 177, 179, 181, 179, 181, 182, 183, 176, 181, 177, 173, 172, 154, 142, 121, 98, 75, 66, 60, 67, 66, 60, 163, 137, 104, 102, 70, 86, 154, 213, 227, 229, 230, 230, 228, 229, 230, 230, 230, 230, 229, 228, 229, 229, 229, 228, 227, 228, 229, 229, 227, 225, 220, 219, 224, 227, 226, 225, 226, 226, 226, 227, 224, 224, 222, 222, 224, 220, 224, 223, 216, 214, 230, 229, 226, 229, 129, 225, 233, 232, 234, 234, 236, 237, 234, 223, 176, 86, 81, 86, 120, 120, 118, 110, 134, 140, 139, 135, 139, 149, 152, 133, 77, 73, 73, 75, 75, 86, 118, 189, 222, 224, 225, 224, 222, 220, 220, 220, 211, 197, 106, 94, 132, 203, 143, 171, 180, 217, 230, 231, 228, 228, 226, 215, 205, 221, 231, 231, 235, 232, 224, 214, 144, 178, 165, 129, 82, 71, 84, 82, 95, 149, 163, 179, 185, 181, 187, 183, 157, 172, 126, 158, 113, 120, 226, 230, 231, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 230, 231, 232, 232, 232, 231, 231, 232, 232, 232, 232, 232, 232, 233, 234, 233, 233, 233, 234, 235, 236, 235, 233, 230, 214, 189, 187, 176, 178, 182, 181, 176, 176, 185, 183, 177, 166, 155, 138, 125, 109, 140, 152, 64, 55, 87, 98, 94, 89, 84, 83, 76, 78, 77, 95, 112, 124, 139, 150, 159, 163, 162, 166, 166, 168, 170, 165, 161, 147, 140, 121, 101, 84, 74, 70, 67, 70, 74, 89, 115, 126, 139, 153, 102, 128, 110, 73, 96, 172, 216, 228, 230, 231, 229, 229, 230, 230, 230, 231, 229, 228, 229, 229, 230, 228, 228, 227, 227, 227, 226, 224, 222, 220, 223, 225, 227, 225, 224, 227, 224, 225, 226, 224, 225, 223, 225, 224, 224, 221, 217, 212, 231, 227, 229, 230, 134, 228, 234, 233, 234, 235, 236, 238, 235, 224, 181, 85, 79, 82, 111, 107, 78, 76, 100, 124, 131, 140, 140, 143, 144, 103, 69, 68, 74, 74, 75, 81, 101, 186, 217, 222, 220, 221, 218, 212, 218, 220, 207, 199, 109, 90, 136, 200, 158, 172, 185, 217, 230, 228, 228, 229, 228, 227, 219, 222, 229, 228, 232, 231, 227, 216, 175, 189, 192, 175, 107, 78, 85, 86, 105, 160, 155, 169, 180, 184, 184, 178, 156, 166, 125, 154, 107, 128, 226, 229, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 231, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 232, 232, 233, 232, 232, 232, 234, 233, 234, 233, 234, 234, 235, 236, 235, 235, 235, 232, 222, 191, 177, 148, 168, 180, 185, 177, 180, 182, 185, 185, 178, 161, 143, 122, 192, 94, 55, 63, 87, 87, 84, 80, 78, 73, 66, 67, 63, 70, 61, 63, 76, 79, 90, 100, 107, 108, 110, 113, 107, 94, 89, 76, 63, 51, 66, 70, 74, 86, 106, 129, 153, 180, 202, 200, 173, 148, 135, 88, 131, 99, 75, 105, 184, 221, 229, 230, 229, 228, 229, 228, 230, 230, 228, 228, 228, 229, 229, 227, 229, 227, 227, 228, 227, 224, 222, 221, 223, 225, 226, 226, 226, 225, 221, 224, 224, 223, 224, 223, 224, 224, 219, 219, 218, 214, 233, 230, 230, 231, 144, 229, 234, 233, 235, 236, 237, 238, 235, 222, 175, 80, 85, 76, 96, 97, 81, 86, 80, 94, 117, 128, 138, 144, 136, 84, 74, 66, 70, 70, 70, 77, 85, 173, 209, 210, 210, 209, 207, 200, 202, 199, 184, 180, 108, 87, 135, 204, 153, 168, 182, 208, 230, 228, 228, 229, 228, 229, 229, 228, 229, 231, 232, 231, 227, 211, 166, 152, 154, 175, 147, 88, 95, 96, 118, 161, 161, 167, 173, 172, 173, 160, 139, 171, 126, 152, 109, 130, 227, 229, 230, 230, 230, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 231, 232, 233, 232, 232, 232, 234, 233, 234, 233, 232, 234, 235, 236, 235, 235, 236, 236, 234, 226, 198, 147, 126, 159, 181, 180, 179, 179, 178, 185, 180, 170, 132, 138, 162, 69, 59, 73, 99, 95, 90, 89, 93, 84, 75, 67, 69, 62, 54, 53, 55, 55, 52, 54, 55, 57, 57, 52, 56, 47, 44, 50, 56, 69, 74, 102, 155, 175, 191, 202, 213, 223, 227, 228, 216, 149, 150, 142, 94, 145, 85, 69, 118, 195, 224, 229, 229, 228, 229, 229, 230, 231, 228, 227, 228, 229, 229, 228, 227, 226, 227, 227, 226, 225, 222, 222, 223, 226, 226, 225, 227, 224, 223, 223, 224, 224, 223, 224, 222, 223, 221, 221, 219, 212, 232, 230, 228, 230, 130, 224, 233, 235, 235, 236, 236, 235, 234, 223, 169, 78, 78, 73, 79, 84, 124, 117, 99, 150, 192, 157, 160, 170, 155, 87, 92, 99, 103, 96, 88, 93, 98, 139, 164, 154, 145, 134, 125, 107, 98, 93, 79, 141, 104, 90, 134, 204, 157, 173, 182, 202, 229, 229, 230, 229, 230, 232, 231, 232, 231, 232, 232, 230, 226, 188, 126, 144, 126, 154, 176, 155, 127, 104, 146, 164, 160, 133, 133, 131, 136, 132, 122, 163, 126, 149, 109, 128, 226, 229, 231, 231, 230, 230, 230, 230, 231, 231, 230, 229, 230, 231, 232, 231, 230, 230, 229, 231, 231, 230, 230, 230, 231, 231, 230, 230, 231, 231, 232, 232, 231, 231, 231, 232, 233, 231, 231, 231, 231, 232, 232, 233, 232, 232, 233, 234, 233, 233, 233, 233, 235, 235, 235, 235, 235, 236, 237, 235, 229, 207, 152, 120, 140, 172, 183, 181, 176, 172, 177, 168, 116, 205, 90, 57, 65, 79, 104, 98, 94, 89, 87, 80, 76, 77, 75, 72, 73, 73, 73, 76, 73, 66, 65, 68, 75, 77, 83, 67, 77, 75, 69, 78, 117, 193, 216, 222, 228, 228, 230, 232, 234, 232, 225, 202, 106, 65, 54, 131, 135, 68, 72, 144, 210, 227, 229, 228, 229, 230, 230, 230, 229, 228, 228, 228, 228, 227, 225, 225, 225, 225, 227, 224, 223, 221, 226, 226, 226, 226, 226, 225, 224, 223, 223, 224, 224, 222, 222, 222, 221, 223, 220, 212, 233, 229, 228, 229, 128, 222, 233, 234, 234, 235, 236, 235, 232, 221, 159, 81, 78, 77, 109, 131, 180, 149, 173, 178, 214, 203, 208, 197, 177, 104, 126, 132, 150, 92, 89, 91, 86, 83, 93, 93, 92, 87, 85, 81, 78, 78, 77, 129, 94, 92, 129, 195, 163, 172, 182, 204, 228, 230, 230, 229, 230, 231, 232, 230, 229, 230, 231, 231, 229, 214, 187, 184, 175, 200, 196, 183, 166, 127, 178, 182, 166, 150, 146, 151, 160, 154, 143, 164, 131, 154, 113, 126, 226, 229, 231, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 230, 230, 229, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 231, 232, 232, 232, 232, 231, 233, 234, 233, 233, 233, 234, 234, 235, 235, 235, 235, 236, 237, 237, 236, 231, 220, 171, 117, 121, 156, 176, 179, 176, 169, 135, 166, 141, 61, 65, 66, 112, 133, 121, 110, 95, 85, 82, 72, 75, 75, 69, 74, 69, 72, 74, 85, 95, 97, 96, 92, 78, 88, 91, 79, 72, 87, 152, 210, 228, 229, 231, 232, 230, 229, 232, 232, 233, 231, 223, 193, 93, 54, 67, 158, 122, 70, 90, 181, 223, 229, 228, 230, 230, 229, 230, 229, 227, 228, 229, 229, 228, 227, 226, 228, 228, 227, 226, 224, 224, 227, 227, 225, 227, 227, 224, 227, 224, 223, 224, 221, 222, 221, 220, 216, 216, 210, 204, 233, 229, 228, 229, 127, 224, 232, 235, 235, 233, 235, 234, 231, 220, 164, 77, 74, 88, 138, 166, 198, 172, 188, 181, 213, 213, 215, 200, 173, 113, 125, 148, 127, 84, 78, 77, 81, 85, 89, 88, 92, 91, 85, 80, 82, 75, 80, 152, 100, 92, 148, 200, 157, 171, 187, 205, 230, 231, 230, 230, 230, 231, 230, 230, 230, 230, 230, 231, 229, 218, 176, 175, 178, 191, 189, 176, 174, 184, 203, 194, 172, 157, 161, 160, 167, 161, 143, 176, 134, 163, 113, 123, 225, 230, 230, 230, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 229, 229, 231, 231, 231, 230, 230, 230, 232, 232, 231, 230, 231, 232, 232, 232, 231, 230, 231, 232, 233, 232, 231, 232, 233, 234, 233, 231, 232, 233, 234, 233, 232, 233, 234, 235, 237, 237, 237, 236, 233, 226, 192, 127, 108, 127, 157, 170, 178, 138, 209, 84, 48, 53, 74, 134, 144, 141, 139, 125, 125, 111, 103, 103, 97, 98, 101, 106, 118, 120, 118, 107, 97, 87, 90, 90, 85, 76, 78, 105, 181, 220, 229, 230, 230, 230, 231, 231, 229, 230, 231, 233, 234, 231, 220, 194, 91, 58, 108, 172, 124, 70, 125, 206, 227, 228, 229, 230, 229, 230, 230, 228, 229, 229, 227, 229, 228, 228, 229, 229, 228, 228, 226, 226, 225, 228, 226, 223, 222, 219, 218, 208, 203, 198, 189, 187, 176, 171, 162, 153, 143, 137, 233, 229, 229, 228, 132, 224, 233, 234, 235, 234, 234, 234, 230, 222, 162, 80, 77, 85, 154, 172, 195, 182, 186, 188, 212, 215, 215, 203, 179, 115, 130, 154, 81, 64, 72, 82, 84, 88, 90, 90, 92, 90, 86, 78, 65, 57, 61, 143, 102, 94, 144, 200, 165, 174, 190, 205, 230, 232, 230, 230, 229, 231, 231, 231, 229, 229, 229, 232, 229, 217, 181, 162, 157, 166, 168, 146, 178, 216, 209, 200, 177, 161, 155, 158, 161, 160, 144, 170, 134, 164, 114, 120, 224, 229, 231, 231, 231, 229, 229, 230, 231, 230, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 230, 231, 232, 232, 232, 231, 231, 231, 232, 232, 231, 230, 231, 232, 232, 233, 231, 231, 233, 234, 233, 232, 233, 232, 233, 233, 231, 233, 234, 236, 236, 237, 236, 237, 238, 237, 232, 211, 151, 105, 96, 123, 135, 185, 171, 40, 36, 42, 92, 130, 135, 142, 146, 145, 146, 138, 136, 136, 131, 131, 129, 123, 120, 106, 95, 96, 99, 98, 83, 74, 72, 98, 158, 199, 225, 230, 229, 230, 230, 231, 231, 230, 229, 230, 231, 231, 233, 233, 228, 220, 193, 92, 62, 163, 182, 124, 74, 161, 216, 227, 229, 228, 228, 229, 228, 228, 227, 226, 222, 222, 219, 215, 216, 206, 201, 200, 191, 185, 174, 172, 166, 160, 153, 141, 142, 133, 131, 126, 129, 128, 128, 116, 106, 98, 71, 59, 232, 228, 228, 228, 144, 226, 233, 234, 234, 234, 234, 233, 231, 223, 159, 93, 89, 98, 158, 172, 185, 190, 178, 190, 201, 215, 212, 201, 197, 118, 121, 143, 71, 66, 74, 85, 74, 99, 97, 95, 93, 93, 86, 56, 54, 50, 50, 136, 107, 100, 151, 206, 158, 178, 200, 206, 231, 231, 230, 230, 230, 231, 232, 232, 231, 230, 229, 232, 229, 220, 196, 156, 156, 153, 150, 166, 220, 230, 218, 208, 193, 165, 139, 133, 138, 144, 147, 165, 133, 162, 111, 122, 224, 230, 231, 231, 230, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 230, 230, 230, 232, 232, 231, 231, 231, 231, 232, 231, 231, 231, 230, 232, 233, 232, 231, 231, 232, 233, 233, 232, 232, 232, 234, 234, 234, 233, 234, 234, 236, 236, 236, 236, 237, 239, 239, 235, 225, 189, 131, 112, 140, 209, 76, 40, 39, 46, 109, 137, 136, 126, 125, 124, 119, 114, 117, 114, 104, 102, 98, 99, 96, 109, 102, 93, 84, 57, 56, 77, 122, 184, 212, 223, 226, 226, 227, 227, 227, 227, 229, 227, 226, 225, 226, 228, 229, 230, 230, 224, 215, 189, 72, 136, 198, 158, 99, 107, 177, 197, 194, 190, 185, 179, 177, 169, 161, 162, 154, 144, 144, 134, 135, 131, 126, 126, 126, 118, 117, 121, 122, 124, 123, 117, 122, 113, 101, 89, 79, 64, 55, 46, 42, 43, 53, 52, 233, 229, 229, 230, 135, 226, 233, 234, 234, 234, 234, 235, 230, 222, 155, 92, 91, 88, 159, 165, 176, 201, 177, 191, 189, 214, 211, 207, 199, 131, 148, 105, 67, 72, 72, 76, 87, 99, 98, 96, 96, 87, 62, 44, 48, 51, 48, 132, 100, 102, 152, 200, 158, 181, 199, 208, 230, 230, 230, 230, 229, 231, 232, 232, 231, 229, 229, 228, 227, 222, 206, 180, 167, 157, 185, 222, 232, 232, 230, 213, 205, 180, 157, 159, 157, 155, 164, 160, 134, 163, 111, 120, 225, 230, 231, 231, 230, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 232, 231, 231, 230, 230, 231, 231, 232, 231, 230, 230, 232, 232, 232, 231, 231, 231, 232, 232, 231, 231, 231, 232, 233, 232, 231, 231, 232, 233, 233, 232, 231, 232, 233, 234, 234, 233, 233, 234, 235, 236, 235, 236, 237, 238, 239, 240, 237, 235, 226, 187, 185, 175, 50, 34, 35, 46, 106, 137, 141, 138, 140, 147, 139, 136, 131, 111, 124, 109, 121, 112, 100, 89, 57, 45, 39, 38, 40, 52, 64, 91, 114, 125, 137, 148, 153, 156, 157, 155, 155, 153, 147, 154, 152, 153, 148, 155, 153, 148, 127, 109, 68, 80, 94, 89, 94, 95, 107, 112, 110, 115, 109, 119, 106, 106, 108, 113, 120, 115, 116, 118, 116, 118, 112, 113, 116, 117, 112, 102, 88, 79, 74, 60, 54, 43, 41, 42, 44, 50, 67, 79, 94, 100, 106, 112, 233, 230, 230, 232, 147, 227, 234, 232, 233, 234, 235, 235, 231, 221, 143, 78, 75, 89, 159, 164, 175, 198, 176, 193, 185, 214, 211, 203, 203, 136, 159, 74, 65, 74, 68, 77, 93, 99, 95, 103, 94, 81, 47, 46, 46, 45, 47, 138, 103, 96, 147, 197, 156, 189, 205, 212, 230, 230, 230, 229, 230, 230, 231, 230, 229, 229, 229, 229, 230, 225, 215, 219, 219, 212, 225, 230, 232, 233, 233, 226, 216, 197, 165, 152, 157, 147, 155, 160, 134, 170, 113, 135, 227, 230, 231, 232, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 230, 229, 230, 230, 231, 231, 231, 230, 230, 231, 232, 231, 230, 231, 231, 232, 232, 232, 231, 231, 232, 232, 232, 232, 232, 232, 233, 232, 232, 231, 232, 232, 233, 233, 232, 232, 232, 233, 234, 234, 233, 234, 234, 235, 236, 234, 236, 236, 239, 238, 239, 237, 238, 236, 184, 222, 112, 170, 136, 79, 46, 43, 56, 69, 85, 91, 110, 109, 107, 98, 89, 95, 66, 65, 52, 48, 50, 49, 52, 50, 48, 49, 50, 54, 56, 59, 59, 67, 68, 78, 74, 74, 78, 77, 79, 76, 72, 73, 75, 77, 78, 78, 73, 67, 64, 60, 62, 71, 72, 72, 73, 77, 82, 86, 91, 97, 102, 105, 106, 103, 101, 105, 107, 100, 96, 87, 85, 69, 63, 56, 48, 46, 43, 51, 45, 43, 49, 60, 73, 77, 90, 100, 116, 121, 125, 130, 128, 124, 117, 233, 229, 229, 232, 154, 229, 234, 233, 235, 235, 236, 236, 232, 221, 138, 79, 75, 85, 153, 156, 165, 181, 165, 175, 167, 199, 188, 183, 183, 135, 139, 70, 66, 70, 78, 77, 95, 97, 98, 106, 97, 67, 47, 42, 44, 49, 45, 145, 105, 97, 161, 205, 166, 189, 195, 211, 230, 231, 229, 229, 230, 231, 230, 230, 229, 230, 230, 228, 228, 219, 211, 219, 214, 210, 215, 215, 231, 233, 233, 231, 224, 209, 184, 163, 164, 156, 154, 156, 133, 174, 118, 132, 226, 230, 232, 231, 230, 230, 230, 230, 230, 231, 231, 230, 230, 231, 231, 230, 230, 230, 230, 232, 231, 231, 230, 230, 231, 231, 232, 231, 231, 231, 232, 232, 231, 231, 231, 232, 233, 232, 232, 232, 232, 234, 233, 232, 230, 219, 218, 231, 233, 230, 232, 233, 234, 234, 235, 234, 234, 234, 235, 233, 231, 229, 225, 224, 216, 206, 200, 191, 187, 196, 163, 77, 113, 99, 64, 44, 47, 49, 52, 53, 55, 57, 59, 54, 52, 50, 51, 51, 52, 48, 51, 55, 51, 57, 53, 54, 48, 53, 49, 51, 52, 52, 60, 56, 62, 60, 57, 57, 63, 57, 59, 58, 59, 64, 58, 60, 58, 53, 53, 59, 60, 58, 64, 66, 75, 74, 77, 74, 78, 76, 76, 73, 79, 70, 62, 58, 51, 48, 44, 46, 44, 46, 48, 48, 51, 57, 61, 82, 81, 88, 98, 109, 106, 109, 111, 121, 119, 129, 128, 132, 131, 118, 110, 98, 234, 232, 230, 234, 147, 232, 236, 237, 236, 238, 239, 239, 235, 225, 137, 82, 74, 83, 99, 91, 100, 94, 93, 99, 116, 131, 122, 114, 121, 144, 94, 77, 90, 91, 79, 82, 78, 65, 72, 109, 101, 57, 50, 52, 57, 53, 50, 146, 107, 106, 168, 211, 160, 190, 196, 208, 230, 231, 230, 228, 230, 231, 230, 230, 229, 229, 230, 229, 229, 211, 200, 210, 199, 208, 209, 205, 222, 232, 233, 233, 229, 220, 208, 186, 190, 180, 154, 149, 135, 178, 113, 139, 227, 230, 232, 232, 231, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 231, 231, 230, 231, 232, 232, 231, 231, 231, 231, 232, 233, 231, 232, 232, 233, 233, 233, 232, 232, 234, 234, 234, 233, 234, 235, 237, 237, 232, 226, 212, 136, 195, 194, 174, 202, 211, 214, 211, 210, 203, 192, 189, 182, 164, 151, 133, 124, 112, 98, 89, 80, 80, 90, 156, 66, 60, 54, 50, 53, 49, 55, 54, 55, 55, 58, 57, 51, 54, 50, 57, 55, 58, 54, 56, 53, 58, 56, 53, 57, 45, 53, 50, 49, 51, 50, 53, 48, 53, 59, 57, 54, 53, 49, 54, 52, 55, 55, 58, 55, 53, 53, 50, 58, 64, 94, 94, 84, 68, 69, 72, 66, 53, 51, 49, 45, 41, 38, 40, 41, 49, 61, 75, 73, 80, 93, 100, 111, 104, 116, 117, 118, 120, 129, 130, 132, 130, 130, 129, 119, 123, 117, 120, 115, 122, 121, 110, 104, 101, 235, 232, 230, 235, 139, 231, 237, 237, 236, 239, 240, 240, 235, 226, 133, 90, 73, 77, 64, 65, 66, 66, 71, 74, 95, 99, 119, 140, 153, 158, 71, 78, 94, 82, 68, 63, 52, 54, 52, 91, 103, 56, 72, 97, 103, 70, 51, 140, 98, 107, 168, 207, 157, 184, 189, 215, 231, 230, 230, 228, 231, 231, 231, 230, 230, 231, 230, 230, 228, 218, 205, 201, 196, 196, 201, 199, 213, 232, 233, 233, 231, 228, 221, 220, 225, 216, 173, 143, 137, 178, 109, 138, 226, 230, 232, 233, 231, 230, 230, 231, 231, 232, 231, 231, 231, 232, 233, 232, 231, 231, 231, 233, 232, 232, 232, 232, 231, 234, 234, 233, 233, 234, 235, 235, 235, 234, 235, 236, 237, 238, 237, 238, 240, 242, 244, 240, 234, 222, 114, 85, 79, 86, 86, 82, 80, 84, 89, 86, 84, 86, 78, 79, 75, 72, 67, 70, 66, 69, 64, 67, 62, 66, 55, 56, 58, 58, 64, 64, 62, 63, 91, 95, 60, 51, 51, 53, 47, 56, 51, 50, 53, 51, 81, 62, 77, 54, 63, 54, 59, 53, 53, 52, 51, 51, 53, 54, 82, 64, 67, 57, 51, 52, 47, 55, 49, 52, 50, 49, 52, 46, 57, 76, 128, 85, 72, 53, 47, 41, 40, 40, 35, 50, 58, 67, 81, 96, 96, 116, 127, 131, 132, 136, 149, 142, 145, 138, 137, 131, 127, 121, 128, 127, 119, 122, 124, 123, 115, 115, 115, 107, 109, 113, 115, 106, 111, 108, 234, 231, 230, 235, 135, 230, 237, 237, 238, 238, 240, 239, 235, 226, 126, 95, 78, 77, 55, 60, 64, 68, 71, 85, 109, 165, 210, 220, 216, 167, 77, 77, 71, 68, 60, 53, 53, 54, 51, 74, 121, 64, 99, 120, 119, 80, 58, 135, 99, 106, 171, 211, 152, 188, 191, 216, 231, 231, 230, 230, 230, 230, 231, 230, 230, 231, 231, 231, 229, 222, 214, 196, 186, 191, 192, 185, 205, 232, 233, 234, 232, 232, 227, 225, 226, 219, 168, 146, 132, 176, 109, 136, 225, 230, 232, 232, 232, 231, 231, 232, 232, 233, 231, 232, 231, 232, 233, 232, 231, 231, 232, 232, 233, 232, 232, 232, 228, 233, 235, 233, 233, 234, 234, 235, 235, 235, 235, 237, 238, 238, 239, 240, 241, 244, 245, 241, 232, 214, 85, 72, 64, 65, 64, 61, 60, 62, 58, 84, 71, 75, 56, 59, 54, 58, 57, 57, 51, 53, 72, 54, 60, 53, 48, 50, 48, 48, 52, 56, 58, 78, 102, 106, 55, 53, 49, 48, 49, 48, 46, 51, 49, 47, 104, 67, 69, 50, 50, 49, 45, 50, 50, 48, 51, 49, 54, 70, 111, 80, 62, 48, 48, 46, 52, 54, 52, 50, 50, 49, 44, 46, 56, 65, 98, 64, 85, 102, 91, 82, 81, 82, 95, 101, 119, 135, 144, 148, 144, 153, 145, 141, 131, 126, 129, 129, 127, 129, 127, 121, 126, 124, 124, 120, 118, 122, 115, 117, 110, 110, 102, 104, 109, 117, 125, 131, 122, 117, 233, 232, 229, 234, 144, 231, 237, 237, 236, 238, 240, 238, 234, 224, 121, 87, 76, 81, 63, 70, 86, 103, 86, 135, 186, 227, 231, 231, 220, 123, 60, 73, 59, 84, 80, 56, 60, 73, 65, 68, 128, 73, 88, 110, 114, 87, 64, 139, 97, 102, 170, 210, 152, 185, 180, 216, 230, 231, 229, 229, 230, 231, 230, 231, 229, 231, 232, 231, 229, 219, 211, 188, 185, 186, 183, 163, 202, 232, 233, 233, 232, 232, 231, 226, 225, 219, 169, 145, 132, 167, 113, 137, 227, 230, 232, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 232, 233, 232, 230, 231, 232, 232, 233, 232, 232, 232, 230, 233, 234, 233, 233, 234, 234, 230, 233, 234, 236, 238, 239, 239, 240, 241, 242, 244, 245, 241, 232, 206, 85, 68, 57, 59, 51, 60, 60, 60, 50, 90, 82, 61, 63, 50, 44, 50, 51, 50, 49, 47, 83, 56, 58, 53, 48, 46, 45, 44, 48, 48, 56, 96, 102, 111, 51, 48, 45, 45, 46, 47, 46, 50, 45, 46, 98, 67, 68, 47, 50, 45, 43, 49, 46, 46, 54, 47, 52, 82, 106, 83, 60, 48, 47, 45, 46, 49, 47, 51, 43, 48, 47, 46, 68, 65, 74, 66, 109, 121, 122, 127, 138, 137, 145, 149, 149, 144, 131, 124, 120, 121, 116, 122, 122, 126, 138, 129, 122, 121, 113, 112, 111, 117, 114, 122, 119, 117, 123, 121, 116, 119, 118, 114, 113, 119, 112, 112, 102, 90, 233, 230, 229, 233, 135, 231, 236, 236, 235, 236, 238, 236, 231, 220, 115, 85, 74, 93, 90, 122, 162, 152, 111, 160, 225, 233, 236, 229, 217, 89, 59, 77, 70, 86, 74, 60, 72, 100, 81, 82, 138, 101, 74, 95, 84, 81, 62, 139, 92, 108, 168, 203, 154, 186, 186, 218, 230, 230, 230, 230, 230, 230, 229, 227, 229, 229, 231, 231, 228, 212, 206, 190, 189, 189, 179, 175, 224, 233, 233, 233, 233, 232, 232, 228, 227, 220, 169, 145, 131, 157, 106, 142, 228, 231, 231, 232, 232, 231, 231, 232, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 232, 232, 233, 232, 232, 232, 234, 234, 234, 233, 232, 232, 221, 220, 229, 231, 236, 238, 239, 240, 240, 241, 242, 245, 246, 242, 231, 206, 80, 64, 55, 49, 49, 50, 51, 56, 54, 87, 78, 56, 54, 49, 46, 44, 47, 50, 52, 45, 93, 57, 59, 50, 46, 46, 41, 42, 45, 50, 56, 117, 103, 90, 50, 45, 50, 47, 45, 46, 48, 46, 50, 46, 103, 57, 67, 48, 45, 46, 44, 48, 47, 45, 46, 44, 53, 82, 95, 92, 55, 49, 49, 44, 48, 43, 42, 47, 48, 50, 44, 41, 70, 74, 63, 97, 149, 147, 134, 124, 111, 110, 108, 114, 115, 109, 119, 114, 112, 110, 119, 120, 124, 129, 123, 126, 118, 123, 112, 106, 112, 113, 120, 122, 115, 119, 114, 112, 112, 113, 106, 103, 97, 101, 93, 89, 85, 82, 232, 229, 229, 232, 149, 231, 235, 235, 235, 237, 238, 236, 230, 220, 113, 86, 80, 104, 150, 161, 146, 122, 106, 178, 231, 238, 235, 226, 202, 72, 62, 67, 70, 61, 54, 67, 81, 94, 82, 98, 138, 113, 104, 85, 86, 70, 62, 141, 85, 118, 158, 177, 155, 190, 179, 216, 230, 230, 230, 230, 229, 230, 229, 229, 230, 231, 230, 228, 227, 195, 199, 188, 188, 185, 180, 215, 230, 232, 233, 233, 232, 232, 232, 227, 227, 220, 197, 147, 131, 177, 108, 142, 228, 231, 232, 232, 231, 231, 231, 232, 233, 232, 232, 231, 231, 232, 232, 232, 230, 231, 232, 233, 233, 233, 233, 232, 234, 234, 227, 232, 234, 231, 232, 236, 231, 234, 232, 238, 239, 240, 240, 236, 243, 245, 246, 243, 230, 201, 71, 56, 56, 62, 53, 51, 52, 53, 50, 98, 76, 48, 46, 52, 46, 47, 46, 49, 51, 46, 73, 56, 56, 49, 45, 48, 44, 42, 48, 49, 50, 91, 91, 80, 49, 46, 48, 42, 46, 46, 48, 47, 53, 45, 113, 71, 72, 70, 46, 46, 48, 50, 48, 40, 47, 47, 60, 108, 94, 107, 61, 51, 45, 43, 46, 52, 45, 46, 53, 47, 48, 53, 85, 83, 57, 90, 110, 103, 97, 95, 103, 97, 101, 106, 107, 112, 110, 114, 115, 116, 122, 112, 113, 124, 123, 122, 121, 114, 112, 112, 110, 114, 116, 112, 109, 109, 112, 106, 104, 100, 89, 81, 80, 92, 83, 91, 87, 83, 233, 230, 230, 233, 137, 230, 234, 235, 235, 236, 237, 235, 230, 220, 105, 86, 81, 111, 146, 149, 135, 115, 163, 214, 232, 237, 237, 227, 205, 75, 60, 59, 58, 75, 56, 60, 82, 73, 77, 99, 138, 97, 107, 87, 118, 91, 60, 135, 80, 124, 169, 182, 149, 187, 167, 219, 229, 230, 229, 229, 230, 230, 230, 229, 229, 230, 231, 228, 227, 204, 192, 185, 184, 183, 188, 227, 231, 232, 233, 233, 231, 232, 233, 232, 229, 223, 208, 148, 130, 173, 107, 136, 227, 230, 231, 232, 231, 230, 231, 230, 233, 232, 232, 231, 231, 233, 232, 231, 231, 231, 232, 233, 233, 232, 232, 232, 234, 234, 228, 231, 233, 234, 235, 236, 236, 236, 236, 238, 239, 240, 239, 240, 242, 245, 246, 242, 230, 191, 71, 59, 59, 51, 55, 55, 43, 63, 48, 79, 81, 50, 49, 53, 48, 50, 50, 52, 52, 47, 81, 58, 51, 45, 45, 48, 42, 46, 42, 49, 50, 82, 80, 69, 51, 45, 50, 46, 48, 52, 47, 53, 52, 46, 105, 69, 66, 88, 57, 54, 56, 54, 57, 47, 93, 57, 65, 131, 99, 105, 52, 47, 49, 45, 50, 45, 46, 49, 46, 52, 50, 53, 95, 94, 58, 70, 102, 95, 96, 101, 96, 100, 97, 104, 113, 107, 114, 111, 112, 112, 106, 107, 108, 111, 111, 109, 110, 105, 96, 99, 101, 103, 106, 97, 100, 104, 104, 98, 87, 84, 82, 80, 89, 105, 97, 100, 98, 88, 233, 230, 230, 234, 144, 230, 235, 234, 234, 235, 235, 233, 227, 218, 102, 85, 83, 115, 171, 188, 160, 188, 216, 227, 233, 237, 236, 226, 197, 74, 56, 54, 64, 69, 78, 75, 95, 95, 94, 98, 148, 79, 92, 88, 103, 88, 61, 136, 83, 115, 173, 182, 144, 177, 161, 216, 227, 229, 230, 230, 230, 230, 229, 226, 228, 230, 231, 230, 228, 216, 184, 180, 174, 175, 200, 230, 231, 232, 233, 233, 232, 232, 233, 233, 230, 223, 208, 155, 128, 173, 110, 134, 227, 230, 231, 232, 231, 231, 231, 232, 232, 232, 232, 230, 231, 232, 233, 232, 231, 231, 232, 233, 234, 232, 232, 232, 234, 234, 231, 227, 234, 235, 236, 236, 236, 236, 237, 238, 239, 240, 240, 241, 242, 245, 245, 242, 230, 181, 77, 53, 57, 55, 53, 48, 48, 53, 48, 71, 87, 49, 49, 51, 48, 51, 51, 45, 52, 46, 67, 57, 51, 47, 45, 45, 46, 48, 46, 47, 50, 72, 64, 66, 50, 45, 48, 43, 46, 49, 44, 50, 57, 49, 110, 70, 68, 81, 78, 91, 96, 95, 99, 57, 84, 99, 66, 137, 93, 103, 52, 50, 47, 45, 44, 44, 47, 45, 48, 47, 50, 62, 86, 96, 55, 84, 103, 95, 100, 102, 107, 101, 101, 107, 105, 103, 103, 103, 103, 97, 95, 102, 101, 99, 102, 107, 104, 100, 93, 90, 89, 92, 96, 97, 96, 99, 103, 106, 98, 95, 96, 97, 90, 107, 101, 96, 102, 96, 232, 229, 229, 234, 137, 229, 234, 234, 234, 234, 235, 233, 227, 215, 94, 87, 82, 113, 149, 203, 206, 213, 219, 231, 235, 235, 234, 228, 163, 134, 59, 53, 62, 88, 125, 80, 97, 98, 80, 104, 146, 88, 93, 73, 78, 78, 72, 145, 84, 122, 172, 183, 144, 183, 170, 218, 228, 229, 228, 229, 230, 230, 229, 227, 229, 230, 231, 229, 225, 211, 175, 168, 162, 165, 216, 230, 232, 232, 232, 233, 232, 232, 232, 234, 231, 222, 208, 161, 131, 178, 114, 135, 226, 230, 231, 232, 231, 231, 231, 231, 233, 233, 231, 231, 231, 232, 233, 233, 232, 231, 231, 233, 233, 233, 232, 233, 234, 235, 234, 234, 234, 234, 236, 235, 236, 236, 237, 238, 240, 241, 240, 241, 242, 245, 246, 242, 230, 172, 71, 56, 56, 56, 48, 46, 48, 54, 52, 84, 78, 54, 49, 49, 51, 52, 47, 51, 49, 48, 73, 63, 53, 50, 44, 47, 47, 48, 45, 51, 51, 78, 67, 75, 50, 54, 50, 42, 47, 43, 48, 47, 52, 49, 108, 76, 74, 68, 88, 73, 76, 81, 90, 55, 86, 76, 67, 128, 81, 112, 52, 46, 45, 44, 41, 40, 44, 43, 48, 46, 49, 69, 86, 108, 47, 111, 101, 106, 101, 97, 93, 99, 98, 100, 100, 94, 99, 93, 99, 102, 107, 104, 110, 108, 110, 117, 115, 113, 106, 105, 102, 105, 106, 102, 98, 103, 102, 100, 97, 91, 90, 90, 91, 111, 114, 114, 121, 100, 233, 229, 229, 232, 132, 228, 233, 234, 233, 233, 235, 231, 226, 213, 94, 90, 87, 116, 189, 207, 211, 215, 220, 230, 234, 231, 228, 220, 92, 155, 122, 60, 108, 142, 146, 126, 91, 92, 80, 144, 150, 107, 84, 79, 73, 76, 106, 149, 77, 110, 178, 180, 148, 192, 166, 219, 228, 230, 228, 229, 230, 229, 229, 230, 229, 231, 230, 228, 223, 194, 163, 157, 160, 183, 225, 230, 231, 232, 233, 233, 232, 232, 232, 233, 230, 222, 203, 163, 131, 175, 108, 135, 227, 230, 232, 232, 232, 231, 231, 231, 232, 232, 231, 231, 231, 232, 233, 232, 231, 230, 231, 232, 233, 232, 232, 232, 234, 235, 234, 233, 234, 235, 236, 236, 236, 236, 237, 238, 240, 240, 240, 241, 241, 245, 246, 242, 230, 171, 72, 59, 54, 50, 54, 51, 55, 56, 56, 90, 76, 52, 48, 46, 47, 46, 48, 53, 50, 49, 81, 64, 54, 46, 47, 46, 45, 49, 49, 50, 54, 76, 62, 64, 52, 57, 48, 46, 42, 48, 45, 47, 50, 52, 99, 77, 70, 77, 83, 81, 66, 79, 75, 58, 91, 80, 64, 136, 77, 117, 53, 43, 48, 49, 45, 42, 45, 44, 40, 50, 51, 92, 89, 112, 49, 91, 92, 93, 96, 96, 94, 89, 93, 93, 95, 94, 96, 106, 111, 110, 111, 110, 112, 115, 121, 114, 115, 116, 110, 108, 103, 102, 111, 100, 102, 108, 112, 106, 105, 105, 105, 106, 111, 116, 117, 104, 110, 110, 230, 229, 228, 232, 136, 229, 233, 234, 233, 234, 235, 233, 225, 211, 94, 91, 92, 125, 201, 214, 215, 221, 225, 228, 233, 231, 225, 204, 102, 108, 160, 105, 147, 158, 158, 155, 135, 125, 104, 166, 149, 113, 62, 71, 75, 93, 172, 141, 76, 110, 179, 174, 146, 190, 170, 222, 228, 230, 229, 229, 230, 230, 231, 230, 230, 231, 229, 225, 212, 176, 157, 152, 152, 199, 230, 230, 231, 232, 232, 233, 232, 232, 233, 233, 230, 224, 201, 153, 131, 171, 106, 139, 227, 231, 231, 233, 232, 231, 231, 231, 232, 233, 232, 231, 231, 233, 233, 232, 231, 231, 232, 233, 233, 232, 232, 232, 234, 234, 234, 233, 234, 234, 236, 236, 236, 236, 236, 238, 240, 240, 240, 241, 242, 245, 245, 241, 229, 166, 70, 57, 53, 67, 58, 60, 57, 58, 57, 89, 78, 49, 47, 52, 45, 50, 46, 49, 51, 53, 90, 65, 48, 45, 46, 45, 42, 48, 48, 53, 51, 77, 63, 70, 51, 47, 44, 50, 44, 46, 41, 44, 52, 54, 106, 80, 70, 84, 81, 95, 59, 63, 55, 59, 92, 75, 57, 126, 85, 113, 49, 48, 48, 46, 43, 42, 41, 44, 47, 47, 52, 96, 83, 115, 45, 73, 83, 91, 102, 99, 93, 93, 99, 108, 105, 108, 102, 108, 113, 106, 115, 112, 113, 118, 126, 122, 119, 120, 114, 113, 114, 112, 111, 106, 112, 108, 112, 112, 112, 100, 99, 100, 103, 108, 113, 107, 108, 117, 231, 229, 229, 231, 151, 228, 232, 234, 233, 233, 235, 233, 223, 210, 94, 88, 98, 128, 204, 216, 218, 218, 222, 224, 227, 231, 225, 196, 147, 103, 152, 127, 156, 176, 189, 170, 166, 161, 154, 146, 137, 73, 61, 70, 92, 146, 191, 131, 82, 133, 172, 173, 146, 187, 161, 220, 228, 230, 229, 228, 230, 231, 230, 230, 228, 227, 220, 213, 193, 169, 155, 148, 154, 209, 225, 229, 230, 230, 231, 231, 230, 231, 232, 233, 230, 223, 203, 147, 131, 169, 107, 138, 227, 230, 231, 229, 231, 231, 231, 231, 232, 233, 231, 231, 231, 232, 232, 232, 231, 231, 232, 233, 233, 232, 232, 232, 234, 234, 234, 233, 233, 235, 236, 236, 236, 236, 236, 238, 240, 240, 240, 241, 242, 245, 245, 240, 228, 178, 65, 56, 67, 62, 59, 63, 64, 57, 59, 105, 73, 46, 60, 49, 42, 70, 46, 50, 48, 43, 83, 64, 49, 47, 48, 46, 47, 47, 47, 46, 53, 88, 71, 74, 49, 44, 48, 45, 46, 46, 44, 46, 55, 58, 104, 78, 65, 69, 50, 60, 125, 58, 49, 54, 90, 81, 57, 139, 87, 118, 51, 45, 50, 47, 46, 38, 41, 49, 49, 41, 48, 100, 85, 118, 58, 91, 98, 94, 94, 100, 101, 101, 97, 94, 95, 91, 100, 101, 114, 111, 112, 110, 119, 119, 121, 120, 126, 117, 116, 113, 110, 106, 108, 105, 113, 109, 107, 106, 107, 102, 99, 97, 103, 107, 109, 112, 118, 120, 232, 228, 229, 233, 146, 229, 233, 234, 233, 234, 235, 233, 224, 209, 92, 88, 101, 128, 205, 212, 214, 218, 218, 221, 223, 228, 225, 181, 147, 140, 135, 107, 162, 210, 213, 199, 170, 160, 152, 147, 99, 68, 93, 90, 115, 191, 192, 129, 84, 130, 184, 190, 149, 190, 162, 222, 231, 230, 229, 229, 229, 230, 228, 226, 219, 211, 200, 186, 174, 161, 149, 134, 176, 204, 206, 203, 198, 194, 205, 206, 206, 212, 215, 227, 230, 222, 203, 158, 125, 172, 105, 146, 228, 230, 231, 231, 232, 231, 231, 232, 233, 232, 231, 232, 231, 232, 232, 232, 231, 231, 232, 233, 233, 232, 232, 233, 234, 234, 234, 233, 234, 234, 236, 236, 236, 236, 236, 238, 239, 240, 240, 240, 242, 245, 245, 242, 230, 191, 75, 58, 84, 61, 58, 60, 58, 63, 60, 99, 72, 48, 51, 50, 44, 48, 46, 45, 50, 42, 75, 65, 47, 44, 44, 51, 46, 51, 47, 46, 48, 76, 66, 74, 49, 47, 44, 40, 40, 42, 41, 46, 49, 52, 99, 74, 65, 72, 80, 77, 106, 71, 55, 53, 86, 85, 90, 157, 97, 114, 46, 43, 43, 45, 53, 41, 43, 43, 47, 48, 48, 96, 87, 109, 60, 82, 101, 93, 106, 104, 110, 106, 102, 101, 106, 98, 104, 106, 110, 117, 117, 117, 121, 124, 122, 126, 123, 119, 120, 113, 105, 108, 103, 104, 104, 105, 106, 109, 111, 109, 109, 109, 110, 114, 118, 121, 111, 110, 233, 228, 228, 231, 138, 228, 233, 234, 234, 234, 235, 232, 223, 206, 85, 88, 100, 129, 203, 216, 215, 207, 195, 201, 209, 219, 217, 122, 108, 146, 142, 100, 181, 216, 213, 206, 169, 148, 144, 146, 126, 136, 116, 102, 169, 199, 190, 130, 85, 143, 186, 182, 139, 192, 161, 223, 231, 232, 230, 226, 225, 221, 210, 206, 195, 183, 172, 168, 162, 137, 128, 126, 194, 166, 128, 146, 168, 181, 197, 200, 198, 195, 202, 210, 227, 222, 203, 166, 136, 173, 113, 139, 228, 230, 232, 232, 232, 231, 231, 232, 232, 233, 232, 231, 232, 232, 232, 231, 232, 231, 232, 233, 233, 232, 232, 232, 233, 234, 234, 233, 233, 234, 236, 235, 235, 236, 236, 238, 239, 239, 239, 240, 242, 243, 245, 241, 229, 203, 75, 65, 127, 64, 73, 64, 65, 65, 55, 93, 74, 52, 48, 44, 47, 42, 42, 51, 49, 46, 79, 67, 48, 47, 46, 47, 47, 44, 45, 46, 51, 77, 69, 75, 52, 46, 46, 43, 42, 44, 44, 44, 49, 59, 109, 69, 68, 66, 49, 67, 105, 101, 89, 57, 86, 88, 53, 144, 86, 100, 48, 48, 45, 48, 41, 43, 42, 40, 42, 54, 54, 116, 91, 91, 55, 92, 105, 97, 100, 112, 105, 96, 102, 103, 102, 103, 104, 119, 112, 113, 119, 117, 122, 122, 120, 128, 126, 122, 122, 115, 110, 107, 99, 101, 108, 107, 107, 111, 107, 118, 114, 118, 120, 117, 107, 101, 93, 100, 234, 231, 229, 231, 129, 226, 234, 235, 234, 235, 236, 233, 224, 204, 92, 83, 105, 127, 207, 215, 210, 198, 147, 120, 160, 195, 206, 67, 49, 93, 132, 121, 194, 218, 218, 197, 165, 142, 116, 128, 143, 170, 125, 144, 205, 206, 197, 133, 89, 140, 192, 183, 149, 190, 161, 225, 230, 229, 224, 222, 202, 193, 180, 177, 168, 160, 146, 132, 122, 109, 108, 116, 127, 123, 122, 140, 157, 169, 201, 194, 190, 197, 202, 208, 227, 223, 205, 166, 137, 179, 115, 140, 228, 230, 232, 232, 232, 231, 231, 231, 232, 232, 231, 231, 231, 232, 232, 233, 231, 231, 232, 233, 233, 232, 232, 232, 233, 234, 234, 233, 233, 234, 235, 236, 235, 235, 236, 238, 239, 239, 239, 240, 242, 244, 245, 241, 230, 209, 84, 64, 149, 66, 62, 64, 65, 65, 54, 101, 65, 43, 45, 48, 45, 42, 46, 43, 52, 45, 76, 62, 50, 45, 45, 48, 48, 45, 48, 48, 48, 80, 72, 74, 46, 46, 48, 46, 42, 42, 41, 46, 49, 60, 115, 78, 65, 71, 62, 63, 109, 78, 54, 50, 94, 95, 58, 145, 80, 93, 44, 46, 44, 42, 39, 40, 42, 39, 45, 42, 47, 110, 89, 104, 67, 85, 89, 94, 97, 105, 101, 105, 105, 105, 110, 109, 111, 112, 112, 113, 112, 121, 121, 118, 117, 126, 122, 120, 120, 112, 112, 110, 100, 105, 103, 105, 108, 106, 101, 111, 98, 95, 93, 97, 92, 98, 96, 92, 234, 231, 229, 232, 139, 228, 234, 235, 235, 235, 236, 234, 225, 201, 95, 85, 108, 126, 205, 216, 205, 192, 129, 128, 145, 181, 187, 51, 54, 54, 111, 132, 183, 212, 197, 182, 113, 98, 84, 101, 150, 150, 129, 196, 214, 208, 197, 125, 86, 148, 199, 181, 154, 190, 166, 223, 227, 218, 214, 192, 176, 170, 158, 140, 119, 117, 98, 90, 86, 88, 100, 103, 100, 108, 117, 137, 148, 160, 170, 181, 187, 192, 198, 209, 224, 222, 204, 162, 137, 181, 111, 138, 228, 230, 232, 231, 232, 231, 231, 231, 232, 232, 231, 231, 231, 233, 233, 233, 232, 232, 232, 233, 233, 232, 232, 232, 232, 234, 234, 233, 233, 234, 235, 236, 235, 235, 236, 238, 239, 239, 239, 241, 242, 244, 245, 241, 230, 213, 81, 62, 157, 64, 63, 65, 72, 64, 51, 95, 76, 50, 48, 44, 42, 45, 44, 46, 46, 43, 80, 59, 50, 45, 47, 49, 46, 45, 41, 47, 53, 71, 67, 69, 48, 42, 45, 45, 39, 44, 41, 45, 54, 55, 123, 72, 66, 69, 65, 62, 58, 46, 50, 46, 53, 93, 60, 147, 73, 92, 47, 46, 46, 40, 42, 43, 42, 43, 47, 43, 51, 118, 96, 102, 69, 79, 85, 90, 98, 98, 105, 111, 107, 108, 109, 108, 111, 109, 113, 119, 111, 103, 113, 110, 115, 117, 110, 112, 116, 112, 107, 110, 106, 101, 101, 96, 103, 100, 90, 90, 88, 97, 92, 104, 106, 104, 106, 104, 234, 231, 228, 231, 120, 225, 235, 235, 235, 236, 237, 235, 225, 204, 89, 88, 106, 121, 194, 193, 169, 160, 122, 119, 132, 153, 170, 67, 80, 81, 78, 129, 155, 122, 105, 104, 87, 75, 85, 121, 158, 148, 152, 217, 217, 211, 195, 125, 92, 143, 201, 174, 156, 196, 170, 216, 222, 216, 194, 150, 128, 114, 100, 98, 93, 87, 80, 84, 89, 107, 103, 117, 108, 110, 128, 141, 153, 163, 175, 180, 185, 189, 197, 207, 227, 223, 205, 165, 128, 181, 109, 134, 227, 230, 231, 231, 232, 231, 230, 231, 232, 232, 231, 231, 231, 232, 233, 233, 232, 232, 232, 233, 233, 233, 232, 233, 233, 234, 234, 233, 233, 234, 235, 236, 236, 236, 236, 237, 239, 240, 240, 241, 242, 244, 245, 242, 232, 219, 82, 53, 121, 60, 66, 63, 62, 62, 47, 89, 57, 47, 42, 45, 48, 45, 49, 47, 56, 42, 82, 61, 55, 45, 44, 45, 41, 43, 43, 48, 49, 77, 72, 73, 50, 47, 49, 41, 43, 39, 45, 51, 49, 49, 114, 70, 64, 71, 64, 59, 70, 60, 78, 48, 85, 48, 51, 129, 72, 91, 51, 43, 43, 47, 41, 41, 40, 41, 47, 44, 46, 94, 95, 89, 81, 88, 88, 91, 97, 106, 109, 115, 121, 116, 113, 108, 111, 115, 112, 113, 109, 105, 109, 111, 108, 113, 113, 112, 107, 98, 94, 90, 94, 96, 102, 96, 105, 95, 97, 93, 95, 97, 109, 108, 114, 116, 106, 102, 234, 232, 231, 233, 150, 230, 235, 237, 236, 238, 239, 237, 227, 207, 91, 84, 100, 108, 167, 102, 80, 96, 103, 107, 119, 137, 160, 110, 82, 59, 60, 132, 144, 84, 91, 97, 83, 74, 105, 130, 151, 136, 183, 216, 213, 203, 194, 115, 92, 145, 179, 144, 155, 199, 180, 218, 217, 206, 172, 153, 157, 170, 171, 172, 166, 145, 131, 129, 135, 142, 146, 152, 152, 135, 142, 147, 167, 187, 185, 185, 184, 187, 189, 207, 226, 224, 209, 171, 129, 176, 106, 141, 228, 230, 231, 231, 232, 231, 231, 231, 232, 232, 231, 231, 230, 232, 232, 233, 232, 232, 232, 233, 234, 233, 232, 233, 234, 234, 234, 233, 233, 234, 235, 236, 236, 236, 236, 238, 239, 240, 240, 241, 242, 244, 246, 242, 234, 220, 82, 51, 67, 73, 67, 80, 64, 56, 48, 91, 56, 47, 50, 49, 44, 47, 45, 47, 48, 47, 80, 61, 54, 47, 45, 45, 46, 50, 45, 43, 49, 70, 73, 75, 48, 47, 45, 42, 42, 45, 41, 48, 47, 48, 119, 70, 62, 73, 56, 62, 89, 91, 90, 56, 87, 61, 54, 124, 82, 90, 53, 46, 43, 48, 41, 40, 38, 43, 46, 47, 52, 83, 100, 97, 66, 97, 124, 122, 118, 108, 103, 98, 101, 99, 98, 93, 92, 101, 100, 111, 108, 98, 106, 110, 113, 117, 114, 109, 102, 96, 91, 95, 98, 99, 102, 105, 107, 102, 104, 105, 104, 108, 108, 110, 112, 108, 98, 85, 235, 232, 231, 233, 136, 229, 237, 238, 238, 239, 240, 238, 228, 206, 92, 81, 97, 105, 145, 78, 87, 86, 98, 107, 104, 116, 107, 45, 41, 44, 46, 131, 147, 95, 67, 73, 96, 90, 143, 157, 173, 181, 208, 220, 213, 198, 189, 107, 92, 157, 190, 143, 144, 201, 163, 218, 219, 195, 157, 170, 193, 196, 203, 203, 206, 189, 162, 167, 168, 170, 178, 175, 173, 173, 160, 170, 165, 186, 177, 164, 167, 174, 192, 204, 225, 227, 220, 176, 125, 185, 109, 141, 228, 231, 231, 231, 232, 231, 231, 231, 232, 232, 232, 232, 231, 231, 232, 232, 232, 232, 232, 234, 234, 233, 232, 232, 233, 234, 234, 234, 234, 235, 235, 236, 236, 236, 237, 238, 239, 240, 240, 241, 242, 244, 246, 243, 236, 225, 95, 57, 55, 63, 56, 60, 62, 52, 46, 93, 59, 51, 46, 41, 42, 50, 41, 45, 50, 47, 74, 59, 55, 51, 48, 52, 50, 46, 47, 46, 52, 58, 73, 77, 50, 49, 48, 43, 39, 44, 46, 48, 46, 44, 108, 64, 70, 84, 58, 69, 52, 51, 62, 44, 71, 85, 65, 104, 79, 80, 49, 42, 43, 42, 44, 39, 40, 43, 40, 46, 51, 80, 98, 108, 56, 112, 130, 117, 115, 105, 100, 93, 96, 96, 98, 103, 97, 102, 106, 112, 105, 111, 105, 110, 112, 108, 112, 109, 100, 107, 97, 103, 105, 105, 103, 107, 107, 105, 94, 95, 93, 90, 103, 101, 99, 110, 104, 94, 235, 231, 232, 234, 143, 231, 237, 238, 239, 239, 239, 237, 228, 201, 90, 78, 97, 88, 117, 82, 99, 91, 86, 82, 89, 108, 80, 37, 38, 48, 47, 141, 164, 134, 103, 116, 143, 176, 209, 210, 195, 197, 209, 218, 213, 202, 186, 111, 102, 164, 201, 140, 155, 209, 174, 220, 220, 182, 182, 166, 189, 189, 196, 197, 204, 190, 164, 163, 168, 175, 170, 177, 176, 177, 175, 158, 163, 145, 148, 168, 166, 174, 186, 200, 225, 227, 222, 186, 126, 178, 109, 136, 228, 231, 231, 231, 231, 231, 231, 231, 232, 233, 232, 231, 231, 232, 233, 233, 232, 232, 232, 234, 233, 232, 233, 232, 233, 234, 235, 234, 234, 234, 236, 236, 236, 236, 237, 238, 240, 239, 240, 241, 242, 244, 246, 244, 238, 227, 111, 48, 52, 44, 52, 57, 53, 43, 43, 102, 62, 52, 47, 44, 47, 46, 45, 47, 49, 48, 67, 55, 56, 46, 41, 41, 42, 47, 46, 44, 48, 58, 74, 76, 51, 47, 48, 46, 42, 40, 42, 50, 42, 45, 103, 62, 75, 87, 62, 62, 53, 61, 52, 47, 69, 66, 55, 97, 83, 87, 46, 43, 47, 41, 45, 39, 42, 42, 44, 42, 51, 64, 94, 100, 50, 94, 89, 100, 101, 96, 103, 103, 100, 103, 104, 99, 99, 99, 98, 108, 105, 108, 106, 108, 112, 111, 113, 111, 110, 107, 104, 107, 99, 97, 98, 106, 107, 103, 98, 95, 92, 93, 105, 100, 102, 114, 107, 98, 234, 232, 232, 235, 158, 232, 237, 238, 238, 239, 239, 237, 228, 198, 90, 74, 87, 75, 88, 85, 97, 102, 85, 98, 87, 112, 61, 32, 38, 42, 45, 152, 167, 164, 154, 142, 158, 172, 202, 216, 194, 203, 211, 220, 218, 202, 187, 104, 99, 162, 206, 145, 153, 207, 156, 217, 217, 166, 178, 143, 160, 167, 166, 171, 182, 184, 153, 160, 161, 162, 164, 167, 165, 166, 166, 155, 153, 143, 144, 155, 157, 170, 179, 197, 221, 227, 224, 202, 131, 184, 110, 142, 229, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 232, 232, 232, 232, 232, 232, 234, 233, 233, 233, 232, 233, 234, 234, 234, 234, 234, 235, 236, 236, 236, 236, 237, 239, 239, 239, 240, 241, 244, 246, 244, 239, 227, 127, 52, 54, 49, 46, 51, 49, 44, 47, 91, 60, 56, 49, 49, 43, 45, 42, 41, 43, 46, 64, 59, 58, 45, 42, 42, 42, 47, 44, 49, 53, 53, 87, 76, 59, 45, 44, 41, 40, 42, 40, 46, 48, 43, 93, 60, 71, 76, 52, 51, 45, 79, 70, 52, 64, 61, 53, 73, 78, 91, 49, 42, 45, 40, 43, 36, 39, 38, 42, 43, 48, 61, 107, 112, 58, 91, 87, 98, 93, 96, 103, 91, 92, 93, 105, 104, 105, 112, 105, 102, 100, 102, 97, 107, 109, 109, 110, 108, 106, 105, 97, 94, 97, 94, 100, 106, 100, 100, 97, 96, 99, 96, 98, 110, 104, 115, 115, 96, 235, 232, 231, 236, 135, 233, 237, 238, 238, 239, 239, 237, 228, 193, 83, 72, 86, 73, 97, 82, 95, 95, 93, 83, 99, 127, 52, 38, 39, 45, 51, 157, 163, 153, 115, 87, 88, 136, 204, 215, 202, 212, 219, 220, 218, 204, 186, 100, 109, 156, 211, 137, 160, 202, 156, 218, 219, 183, 180, 127, 121, 113, 109, 117, 134, 152, 139, 148, 147, 151, 153, 160, 158, 158, 154, 153, 146, 143, 152, 157, 158, 167, 173, 192, 218, 223, 223, 210, 128, 183, 108, 146, 228, 230, 231, 232, 232, 231, 230, 231, 232, 231, 231, 231, 231, 231, 232, 226, 231, 232, 233, 234, 234, 233, 233, 233, 234, 234, 234, 233, 233, 234, 235, 236, 236, 236, 236, 238, 239, 240, 240, 240, 242, 244, 246, 244, 240, 227, 141, 52, 44, 46, 49, 50, 49, 44, 51, 80, 63, 59, 48, 47, 50, 41, 41, 51, 45, 48, 61, 60, 57, 45, 44, 41, 46, 47, 49, 49, 52, 46, 77, 73, 47, 46, 51, 52, 45, 43, 43, 49, 51, 49, 96, 61, 78, 72, 67, 55, 45, 68, 56, 45, 66, 69, 50, 70, 83, 75, 46, 43, 45, 39, 37, 43, 37, 40, 42, 42, 52, 50, 97, 103, 52, 76, 80, 96, 102, 94, 102, 98, 94, 103, 108, 97, 100, 99, 97, 105, 114, 114, 120, 124, 116, 112, 104, 108, 102, 104, 103, 99, 108, 101, 106, 108, 105, 109, 104, 108, 97, 97, 93, 100, 91, 89, 88, 69, 236, 231, 231, 235, 133, 232, 237, 238, 238, 239, 239, 237, 227, 189, 86, 76, 92, 92, 118, 82, 84, 92, 91, 80, 128, 134, 43, 40, 43, 52, 59, 151, 150, 105, 96, 95, 86, 114, 189, 216, 181, 206, 220, 222, 216, 199, 176, 98, 109, 153, 209, 142, 161, 205, 164, 227, 227, 212, 200, 182, 121, 119, 134, 129, 106, 110, 115, 114, 127, 136, 136, 146, 152, 145, 145, 142, 131, 140, 137, 152, 153, 158, 168, 188, 214, 217, 220, 213, 124, 180, 102, 150, 228, 231, 231, 232, 232, 231, 231, 231, 232, 232, 231, 231, 230, 232, 230, 229, 230, 231, 232, 234, 234, 233, 233, 233, 233, 234, 234, 233, 233, 234, 236, 235, 236, 236, 236, 238, 239, 240, 240, 240, 242, 244, 246, 244, 241, 228, 161, 57, 49, 43, 46, 50, 43, 45, 49, 62, 66, 61, 45, 47, 45, 42, 43, 47, 42, 47, 52, 58, 59, 46, 43, 46, 41, 42, 51, 48, 47, 48, 77, 65, 51, 44, 44, 42, 43, 46, 42, 42, 47, 48, 79, 72, 88, 92, 66, 72, 53, 61, 49, 41, 52, 71, 48, 54, 93, 68, 52, 44, 43, 41, 37, 37, 38, 39, 40, 41, 44, 41, 96, 107, 60, 101, 140, 133, 120, 102, 101, 96, 95, 92, 98, 97, 103, 98, 101, 104, 115, 114, 111, 111, 113, 117, 113, 113, 110, 112, 105, 99, 108, 104, 104, 103, 101, 97, 93, 93, 82, 74, 69, 71, 75, 81, 89, 92, 235, 233, 231, 235, 152, 233, 237, 237, 238, 239, 238, 237, 227, 185, 89, 79, 105, 117, 139, 99, 101, 93, 84, 80, 115, 119, 39, 39, 42, 53, 83, 136, 100, 100, 96, 92, 68, 71, 152, 184, 167, 191, 212, 219, 202, 188, 152, 94, 109, 135, 187, 148, 156, 202, 168, 228, 232, 231, 225, 215, 187, 114, 107, 110, 113, 103, 90, 91, 108, 113, 119, 129, 126, 135, 134, 136, 127, 124, 136, 159, 145, 151, 163, 192, 214, 215, 220, 217, 128, 183, 100, 146, 228, 230, 231, 232, 232, 231, 231, 231, 232, 231, 231, 231, 231, 232, 232, 232, 232, 232, 232, 234, 233, 233, 232, 232, 234, 234, 234, 234, 234, 234, 235, 235, 236, 236, 236, 238, 239, 240, 240, 240, 242, 244, 246, 245, 241, 228, 182, 63, 49, 54, 47, 45, 43, 40, 45, 51, 69, 58, 45, 44, 47, 44, 40, 45, 41, 47, 47, 62, 54, 42, 47, 44, 37, 44, 47, 49, 50, 43, 76, 61, 50, 44, 44, 46, 40, 46, 43, 46, 41, 45, 65, 72, 83, 98, 76, 56, 45, 60, 47, 59, 68, 67, 51, 47, 94, 63, 53, 42, 42, 39, 43, 40, 249, 43, 49, 40, 48, 43, 104, 90, 60, 67, 93, 89, 87, 90, 92, 84, 91, 90, 93, 91, 100, 100, 107, 108, 118, 111, 114, 109, 110, 109, 106, 105, 99, 95, 82, 87, 88, 81, 77, 85, 92, 82, 75, 67, 70, 75, 73, 83, 83, 93, 92, 86, 235, 233, 229, 235, 128, 229, 237, 237, 237, 239, 239, 237, 226, 178, 90, 75, 114, 91, 112, 75, 74, 81, 86, 98, 117, 100, 47, 53, 92, 135, 141, 90, 100, 95, 86, 75, 68, 76, 131, 180, 174, 178, 191, 209, 202, 157, 153, 90, 110, 124, 194, 170, 159, 199, 170, 225, 231, 232, 223, 224, 211, 186, 134, 93, 85, 82, 86, 90, 89, 95, 102, 108, 115, 113, 118, 112, 115, 125, 118, 124, 131, 150, 162, 200, 208, 210, 214, 219, 124, 171, 100, 146, 228, 230, 231, 232, 231, 230, 231, 231, 232, 232, 231, 231, 231, 232, 233, 233, 232, 231, 232, 234, 234, 233, 232, 233, 234, 234, 235, 234, 233, 233, 235, 236, 235, 236, 236, 238, 238, 240, 240, 241, 241, 244, 245, 245, 242, 230, 197, 69, 50, 48, 52, 43, 46, 45, 42, 47, 68, 51, 49, 44, 43, 41, 42, 45, 42, 46, 44, 73, 57, 44, 41, 43, 42, 44, 43, 48, 46, 40, 75, 61, 57, 47, 48, 44, 44, 47, 43, 47, 44, 49, 57, 76, 72, 64, 65, 49, 56, 74, 66, 61, 79, 69, 59, 45, 88, 58, 59, 42, 43, 46, 41, 43, 42, 45, 37, 43, 46, 36, 114, 85, 61, 53, 97, 105, 106, 97, 90, 88, 88, 87, 86, 95, 92, 90, 98, 107, 104, 101, 95, 88, 87, 87, 81, 79, 77, 68, 74, 82, 85, 83, 93, 87, 96, 89, 85, 82, 84, 86, 96, 104, 97, 103, 94, 85, 235, 232, 229, 233, 118, 228, 236, 237, 237, 238, 238, 237, 225, 175, 82, 75, 110, 81, 83, 70, 65, 72, 75, 81, 109, 115, 75, 134, 196, 198, 170, 91, 84, 89, 77, 74, 68, 113, 136, 173, 176, 175, 183, 175, 204, 196, 137, 92, 106, 116, 209, 165, 156, 193, 173, 217, 223, 221, 214, 218, 213, 206, 196, 175, 137, 87, 77, 83, 86, 89, 82, 89, 96, 99, 101, 99, 97, 101, 106, 115, 116, 133, 147, 181, 186, 188, 188, 207, 114, 164, 96, 144, 228, 230, 232, 231, 231, 230, 231, 231, 232, 233, 231, 231, 231, 232, 232, 233, 232, 231, 233, 233, 234, 233, 233, 233, 234, 234, 234, 233, 233, 234, 236, 236, 236, 236, 236, 237, 239, 239, 239, 240, 241, 243, 244, 245, 242, 233, 213, 79, 57, 46, 48, 46, 45, 46, 47, 39, 68, 52, 51, 46, 47, 43, 41, 43, 48, 42, 42, 75, 55, 47, 41, 44, 40, 42, 45, 43, 46, 46, 74, 62, 70, 46, 45, 44, 42, 46, 44, 41, 46, 51, 49, 79, 64, 59, 66, 58, 66, 67, 58, 56, 44, 62, 65, 44, 85, 53, 56, 43, 41, 42, 41, 38, 45, 41, 40, 41, 38, 41, 88, 74, 65, 49, 96, 111, 106, 100, 89, 84, 77, 82, 74, 77, 80, 78, 77, 94, 80, 91, 91, 91, 89, 88, 82, 83, 83, 78, 84, 93, 97, 92, 93, 98, 106, 97, 100, 98, 92, 99, 99, 98, 102, 102, 100, 93, 235, 232, 229, 234, 141, 231, 236, 238, 238, 239, 237, 236, 225, 170, 73, 76, 108, 81, 89, 68, 65, 68, 70, 81, 134, 107, 65, 114, 203, 200, 159, 84, 67, 69, 78, 94, 125, 152, 165, 173, 176, 97, 105, 112, 145, 167, 128, 95, 94, 141, 222, 172, 156, 191, 150, 162, 164, 152, 146, 150, 146, 137, 137, 131, 112, 93, 80, 80, 81, 84, 82, 80, 82, 89, 84, 85, 87, 79, 84, 77, 78, 81, 89, 100, 90, 101, 113, 125, 105, 132, 85, 142, 228, 230, 232, 231, 231, 230, 231, 232, 232, 233, 231, 231, 231, 232, 232, 233, 232, 232, 233, 233, 233, 233, 233, 233, 233, 234, 234, 233, 233, 233, 235, 234, 235, 236, 235, 237, 238, 238, 237, 240, 239, 241, 242, 243, 240, 236, 223, 127, 69, 52, 50, 45, 45, 43, 45, 42, 60, 51, 52, 45, 42, 39, 44, 43, 40, 45, 41, 62, 52, 53, 43, 44, 42, 43, 42, 46, 49, 42, 61, 57, 70, 44, 43, 42, 45, 43, 45, 44, 44, 47, 46, 88, 62, 61, 65, 48, 44, 40, 40, 60, 41, 61, 61, 51, 80, 53, 61, 40, 40, 43, 39, 37, 38, 40, 42, 39, 39, 38, 67, 76, 63, 46, 94, 96, 99, 92, 83, 76, 72, 76, 82, 78, 81, 85, 95, 98, 98, 101, 106, 102, 108, 97, 97, 100, 99, 98, 103, 110, 105, 99, 97, 110, 106, 100, 104, 97, 93, 99, 102, 111, 112, 104, 105, 103, 235, 231, 231, 235, 133, 231, 237, 239, 239, 240, 239, 236, 226, 167, 72, 78, 96, 86, 88, 65, 59, 58, 67, 89, 157, 112, 63, 72, 192, 200, 142, 84, 72, 74, 102, 109, 138, 133, 117, 138, 133, 61, 89, 73, 76, 77, 87, 94, 106, 126, 220, 178, 151, 179, 105, 102, 103, 96, 88, 81, 78, 79, 82, 80, 78, 81, 82, 83, 82, 89, 81, 81, 84, 87, 83, 81, 83, 79, 81, 85, 84, 83, 85, 91, 94, 97, 97, 95, 98, 112, 79, 128, 227, 230, 231, 232, 232, 231, 230, 231, 232, 232, 231, 231, 231, 232, 233, 233, 232, 232, 232, 233, 233, 233, 233, 232, 234, 234, 234, 233, 232, 233, 234, 232, 234, 235, 234, 236, 237, 237, 235, 236, 237, 236, 239, 240, 238, 239, 231, 207, 118, 73, 54, 47, 52, 50, 46, 44, 56, 48, 49, 45, 39, 41, 46, 46, 42, 42, 38, 69, 49, 55, 42, 42, 39, 44, 46, 47, 46, 43, 54, 64, 67, 45, 45, 42, 45, 43, 44, 44, 48, 46, 46, 83, 55, 58, 64, 54, 41, 42, 42, 46, 45, 88, 72, 62, 62, 59, 52, 44, 42, 41, 37, 38, 48, 37, 42, 38, 33, 39, 52, 62, 78, 39, 82, 100, 98, 91, 89, 83, 85, 81, 97, 87, 90, 99, 101, 99, 108, 106, 111, 106, 107, 98, 103, 101, 99, 98, 99, 109, 103, 102, 97, 115, 103, 104, 104, 104, 103, 103, 110, 111, 119, 105, 105, 102, 234, 233, 232, 236, 144, 233, 238, 240, 239, 241, 240, 237, 225, 161, 72, 75, 98, 80, 87, 71, 69, 67, 79, 101, 164, 102, 59, 64, 165, 174, 113, 100, 80, 72, 67, 72, 72, 66, 65, 68, 66, 65, 58, 59, 61, 63, 77, 84, 105, 109, 215, 186, 147, 113, 103, 96, 89, 88, 79, 72, 77, 78, 78, 83, 86, 81, 88, 93, 81, 85, 88, 87, 91, 91, 95, 97, 98, 98, 103, 108, 102, 102, 96, 96, 101, 102, 101, 96, 109, 88, 109, 154, 227, 231, 231, 232, 232, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 233, 232, 232, 232, 233, 233, 233, 232, 232, 233, 234, 234, 232, 232, 233, 234, 234, 233, 234, 234, 235, 236, 236, 235, 236, 237, 237, 240, 241, 239, 241, 237, 228, 188, 91, 77, 62, 70, 60, 56, 51, 47, 50, 52, 46, 38, 44, 44, 45, 44, 42, 42, 53, 50, 51, 41, 44, 44, 42, 42, 44, 45, 46, 52, 60, 69, 49, 45, 46, 44, 44, 43, 43, 47, 45, 49, 82, 55, 62, 59, 42, 45, 40, 42, 40, 37, 49, 53, 45, 57, 67, 52, 42, 38, 38, 40, 39, 40, 40, 36, 37, 33, 37, 47, 70, 110, 46, 74, 91, 100, 95, 88, 88, 89, 91, 92, 87, 94, 97, 94, 103, 100, 102, 107, 92, 97, 99, 97, 102, 88, 96, 101, 102, 104, 105, 110, 116, 116, 113, 108, 112, 105, 102, 102, 101, 108, 105, 108, 118, 234, 233, 232, 236, 145, 232, 238, 240, 240, 240, 239, 235, 222, 147, 67, 73, 108, 84, 84, 86, 71, 72, 74, 84, 122, 68, 65, 64, 76, 74, 68, 68, 65, 62, 64, 64, 66, 64, 64, 67, 70, 72, 68, 67, 63, 71, 68, 78, 92, 99, 200, 162, 140, 112, 123, 105, 96, 92, 88, 82, 83, 89, 88, 93, 93, 90, 92, 89, 87, 85, 83, 88, 86, 91, 86, 97, 94, 89, 94, 101, 98, 94, 95, 95, 104, 102, 107, 97, 104, 95, 116, 154, 228, 231, 232, 232, 232, 231, 231, 231, 230, 232, 231, 231, 231, 232, 233, 233, 232, 232, 232, 234, 234, 233, 232, 232, 234, 234, 234, 233, 233, 233, 235, 235, 235, 234, 235, 236, 235, 235, 235, 237, 238, 238, 241, 241, 240, 236, 227, 197, 107, 91, 80, 74, 80, 78, 72, 65, 58, 59, 63, 57, 56, 54, 51, 52, 47, 43, 47, 48, 50, 48, 42, 44, 43, 44, 41, 44, 42, 45, 45, 57, 65, 45, 45, 44, 45, 43, 42, 45, 47, 49, 46, 78, 57, 71, 49, 48, 46, 46, 42, 39, 37, 39, 38, 51, 53, 75, 47, 49, 36, 39, 37, 41, 38, 42, 40, 35, 35, 49, 42, 79, 100, 51, 72, 106, 110, 108, 96, 98, 90, 89, 91, 90, 95, 96, 94, 92, 90, 92, 93, 92, 93, 103, 101, 103, 104, 98, 101, 113, 112, 116, 121, 120, 117, 113, 111, 95, 90, 96, 106, 115, 128, 126, 117, 103, 233, 230, 231, 233, 136, 230, 235, 238, 234, 238, 235, 232, 219, 139, 67, 77, 108, 75, 73, 71, 73, 68, 68, 63, 63, 61, 61, 64, 65, 69, 64, 72, 66, 64, 63, 68, 70, 71, 72, 74, 80, 73, 74, 77, 74, 74, 74, 75, 80, 84, 112, 113, 110, 102, 103, 100, 94, 89, 95, 85, 88, 91, 92, 90, 88, 90, 85, 83, 85, 85, 81, 92, 96, 94, 101, 101, 96, 96, 98, 96, 102, 99, 98, 100, 109, 114, 113, 116, 111, 117, 115, 154, 228, 231, 231, 232, 232, 230, 230, 231, 231, 229, 229, 230, 231, 232, 233, 232, 232, 232, 232, 233, 233, 233, 232, 232, 234, 234, 234, 232, 233, 233, 235, 235, 234, 234, 235, 236, 236, 236, 235, 237, 237, 239, 241, 240, 238, 234, 222, 138, 97, 87, 83, 77, 79, 78, 81, 78, 83, 83, 80, 69, 72, 67, 72, 73, 67, 65, 62, 64, 67, 53, 50, 51, 45, 47, 51, 47, 51, 43, 42, 53, 49, 47, 46, 40, 47, 42, 40, 50, 45, 44, 49, 67, 63, 65, 46, 43, 39, 40, 43, 37, 40, 42, 42, 51, 46, 78, 47, 45, 38, 40, 35, 41, 41, 37, 40, 36, 34, 34, 32, 58, 70, 51, 60, 120, 129, 128, 112, 108, 107, 93, 103, 102, 95, 98, 93, 94, 97, 91, 90, 96, 103, 99, 102, 111, 108, 99, 103, 117, 120, 124, 134, 129, 126, 127, 111, 101, 93, 88, 83, 81, 79, 73, 50, 45, 228, 220, 216, 222, 121, 215, 224, 224, 221, 221, 221, 213, 201, 119, 73, 72, 85, 67, 69, 69, 67, 65, 70, 72, 63, 67, 65, 71, 73, 70, 68, 70, 70, 72, 71, 74, 75, 70, 69, 76, 71, 72, 70, 82, 80, 86, 86, 90, 102, 109, 180, 185, 134, 111, 107, 107, 114, 106, 103, 99, 99, 97, 96, 100, 102, 93, 89, 93, 97, 94, 94, 98, 101, 93, 103, 92, 95, 96, 99, 100, 103, 102, 107, 105, 111, 122, 122, 138, 114, 130, 119, 152, 229, 231, 231, 232, 232, 231, 231, 231, 232, 231, 232, 230, 231, 231, 233, 233, 231, 232, 232, 233, 233, 232, 232, 232, 233, 234, 233, 233, 233, 233, 234, 235, 235, 233, 235, 236, 237, 236, 236, 237, 236, 240, 242, 239, 236, 229, 208, 107, 95, 84, 82, 78, 82, 79, 74, 75, 93, 84, 78, 75, 77, 72, 70, 67, 71, 72, 75, 69, 76, 69, 73, 66, 69, 68, 67, 66, 62, 61, 57, 59, 62, 54, 50, 48, 49, 47, 56, 44, 49, 53, 48, 56, 75, 71, 49, 44, 43, 40, 39, 41, 41, 36, 44, 45, 43, 71, 49, 48, 38, 39, 39, 46, 36, 38, 38, 36, 32, 33, 37, 51, 52, 57, 50, 108, 116, 110, 107, 106, 101, 97, 103, 103, 93, 101, 93, 101, 103, 104, 107, 108, 116, 121, 124, 121, 129, 115, 114, 114, 114, 102, 88, 83, 77, 65, 58, 50, 46, 44, 48, 49, 39, 63, 37, 36, 204, 200, 200, 202, 114, 200, 206, 197, 204, 204, 204, 201, 195, 114, 68, 69, 72, 67, 64, 66, 67, 73, 67, 68, 70, 79, 71, 76, 69, 67, 69, 74, 73, 68, 72, 71, 78, 77, 76, 81, 86, 91, 87, 88, 88, 86, 90, 89, 107, 109, 190, 200, 137, 122, 108, 113, 114, 112, 107, 112, 106, 110, 105, 103, 107, 96, 97, 99, 97, 99, 106, 93, 98, 102, 105, 99, 100, 104, 108, 105, 105, 108, 108, 118, 126, 132, 157, 181, 118, 143, 117, 160, 229, 230, 231, 232, 231, 231, 231, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 232, 232, 233, 233, 232, 232, 232, 233, 234, 234, 233, 233, 233, 234, 235, 235, 234, 235, 236, 237, 236, 236, 237, 237, 240, 240, 240, 236, 227, 200, 106, 89, 86, 79, 80, 81, 83, 82, 76, 96, 88, 89, 76, 73, 71, 75, 77, 71, 71, 74, 78, 85, 78, 69, 74, 69, 74, 73, 75, 74, 73, 77, 70, 75, 76, 65, 65, 58, 69, 66, 62, 62, 63, 67, 81, 100, 96, 69, 57, 54, 46, 40, 47, 44, 41, 43, 45, 41, 62, 49, 52, 39, 39, 43, 37, 37, 40, 39, 37, 37, 37, 49, 48, 61, 54, 44, 98, 126, 120, 115, 108, 111, 103, 107, 109, 96, 104, 105, 109, 107, 105, 103, 95, 100, 95, 87, 85, 74, 66, 59, 58, 61, 50, 44, 44, 43, 39, 40, 36, 38, 37, 38, 50, 45, 45, 44, 54, 207, 209, 205, 208, 105, 207, 208, 214, 212, 210, 211, 207, 201, 108, 72, 73, 73, 69, 68, 68, 68, 68, 65, 66, 67, 69, 74, 74, 72, 79, 78, 74, 79, 71, 80, 77, 80, 81, 82, 89, 88, 89, 82, 93, 94, 92, 88, 93, 104, 123, 188, 179, 140, 173, 128, 140, 142, 141, 137, 141, 137, 138, 133, 129, 114, 100, 102, 100, 102, 100, 102, 103, 112, 104, 105, 110, 112, 116, 113, 122, 122, 130, 137, 163, 170, 178, 196, 209, 134, 158, 125, 156, 229, 231, 232, 231, 231, 231, 230, 231, 231, 232, 230, 231, 232, 232, 233, 233, 231, 232, 232, 233, 233, 233, 232, 232, 233, 234, 233, 232, 233, 233, 234, 235, 234, 234, 234, 236, 236, 236, 235, 235, 237, 240, 238, 238, 235, 225, 192, 98, 98, 89, 81, 81, 83, 86, 84, 76, 105, 86, 85, 76, 75, 74, 75, 72, 78, 79, 78, 85, 93, 80, 74, 75, 76, 71, 72, 75, 74, 78, 69, 84, 76, 77, 73, 73, 68, 78, 78, 73, 72, 68, 75, 79, 91, 73, 64, 64, 62, 55, 51, 52, 56, 48, 56, 51, 44, 53, 48, 50, 42, 39, 37, 36, 39, 42, 45, 40, 41, 43, 42, 48, 57, 53, 55, 73, 108, 95, 86, 65, 68, 71, 67, 72, 70, 64, 58, 59, 58, 50, 53, 50, 46, 50, 47, 43, 50, 41, 43, 45, 40, 43, 49, 48, 47, 48, 50, 44, 50, 49, 54, 54, 55, 56, 54, 55, 205, 208, 208, 208, 121, 208, 211, 215, 214, 213, 210, 210, 199, 134, 80, 67, 69, 76, 72, 71, 68, 71, 73, 71, 73, 76, 75, 76, 83, 82, 81, 78, 78, 75, 82, 86, 84, 83, 90, 92, 96, 94, 98, 104, 107, 114, 106, 92, 107, 124, 195, 171, 146, 190, 156, 180, 181, 175, 177, 181, 177, 169, 160, 138, 114, 100, 103, 103, 105, 109, 109, 114, 119, 117, 120, 123, 117, 119, 125, 128, 131, 145, 146, 168, 180, 185, 209, 212, 132, 159, 127, 162, 229, 230, 232, 231, 231, 231, 230, 231, 232, 232, 231, 231, 231, 232, 232, 233, 231, 232, 232, 233, 233, 233, 232, 232, 234, 233, 233, 233, 233, 233, 233, 234, 233, 233, 233, 235, 236, 236, 234, 235, 236, 239, 238, 237, 234, 224, 184, 96, 91, 90, 91, 87, 85, 86, 83, 84, 104, 85, 85, 76, 76, 82, 78, 81, 83, 87, 77, 91, 92, 82, 77, 74, 73, 78, 79, 76, 80, 74, 84, 90, 89, 83, 79, 78, 73, 80, 70, 77, 71, 72, 70, 81, 101, 100, 80, 74, 74, 69, 73, 68, 67, 64, 68, 69, 62, 55, 55, 50, 46, 44, 44, 37, 45, 44, 45, 47, 43, 46, 55, 65, 75, 88, 107, 88, 75, 57, 59, 42, 42, 44, 44, 51, 46, 41, 41, 42, 40, 42, 43, 45, 41, 43, 47, 47, 48, 52, 51, 59, 70, 70, 77, 72, 74, 74, 67, 62, 64, 66, 68, 66, 72, 62, 60, 60, 199, 206, 205, 209, 120, 206, 209, 212, 213, 210, 208, 207, 197, 115, 87, 84, 82, 83, 83, 74, 77, 78, 81, 85, 83, 87, 83, 84, 94, 96, 84, 84, 78, 82, 82, 91, 99, 102, 112, 132, 126, 99, 117, 129, 151, 152, 127, 103, 121, 123, 173, 201, 156, 197, 160, 185, 189, 187, 188, 181, 175, 145, 127, 116, 110, 109, 112, 107, 107, 115, 117, 114, 126, 129, 128, 129, 129, 130, 135, 146, 143, 145, 148, 172, 180, 188, 211, 209, 128, 158, 121, 160, 229, 231, 232, 232, 231, 230, 231, 231, 231, 232, 231, 231, 232, 232, 232, 233, 232, 231, 232, 233, 233, 233, 232, 232, 234, 234, 233, 233, 233, 233, 233, 234, 233, 233, 234, 234, 236, 237, 233, 235, 236, 239, 237, 236, 233, 224, 179, 104, 94, 96, 87, 86, 84, 82, 84, 81, 111, 87, 87, 81, 78, 80, 71, 81, 84, 80, 80, 92, 88, 88, 83, 79, 79, 76, 79, 81, 77, 84, 76, 91, 88, 83, 75, 75, 72, 75, 79, 80, 74, 71, 81, 78, 102, 88, 80, 75, 72, 70, 74, 66, 69, 77, 76, 76, 68, 70, 68, 69, 66, 63, 61, 53, 58, 55, 58, 54, 53, 51, 70, 88, 117, 134, 132, 139, 93, 73, 60, 41, 46, 44, 50, 44, 51, 52, 56, 58, 50, 55, 53, 55, 59, 66, 67, 57, 63, 60, 64, 75, 72, 74, 80, 85, 86, 90, 83, 77, 80, 81, 83, 94, 98, 99, 99, 102, 202, 204, 204, 210, 130, 207, 209, 210, 214, 212, 208, 203, 195, 113, 85, 88, 83, 91, 90, 84, 85, 87, 79, 83, 96, 81, 90, 94, 121, 121, 104, 98, 92, 89, 99, 110, 120, 130, 137, 148, 142, 140, 147, 156, 169, 144, 129, 96, 122, 132, 158, 195, 159, 188, 157, 189, 191, 191, 184, 176, 147, 116, 122, 126, 123, 119, 116, 116, 121, 123, 127, 129, 130, 130, 135, 136, 129, 132, 138, 149, 147, 149, 154, 170, 181, 186, 208, 202, 126, 159, 123, 158, 228, 229, 231, 232, 231, 231, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 232, 231, 232, 233, 233, 232, 232, 232, 233, 234, 233, 232, 233, 233, 233, 234, 234, 232, 234, 235, 237, 236, 234, 236, 237, 238, 236, 235, 233, 224, 172, 103, 100, 94, 97, 87, 91, 91, 90, 91, 107, 87, 84, 77, 74, 79, 71, 76, 80, 81, 76, 96, 89, 83, 79, 77, 80, 73, 76, 77, 70, 76, 79, 96, 95, 83, 77, 77, 74, 75, 81, 76, 79, 76, 79, 81, 97, 90, 79, 78, 73, 75, 71, 70, 71, 73, 71, 68, 70, 86, 86, 71, 74, 65, 64, 73, 69, 64, 64, 68, 63, 65, 66, 80, 110, 112, 103, 129, 107, 97, 83, 49, 53, 56, 60, 58, 64, 59, 61, 68, 66, 64, 76, 70, 74, 84, 83, 82, 89, 92, 92, 92, 106, 104, 104, 100, 108, 102, 96, 99, 97, 97, 98, 100, 103, 107, 100, 100, 201, 201, 200, 205, 129, 200, 208, 209, 211, 208, 203, 199, 195, 108, 95, 93, 97, 88, 90, 89, 108, 87, 96, 97, 137, 89, 86, 96, 152, 151, 108, 90, 88, 100, 93, 100, 107, 122, 135, 149, 143, 151, 160, 176, 160, 136, 126, 97, 117, 132, 151, 173, 155, 190, 160, 191, 187, 177, 173, 152, 122, 128, 137, 131, 121, 125, 123, 123, 132, 135, 132, 136, 136, 134, 143, 140, 135, 136, 145, 144, 153, 157, 153, 169, 184, 188, 212, 195, 125, 160, 127, 155, 227, 229, 231, 232, 231, 231, 230, 231, 231, 232, 231, 231, 232, 232, 233, 233, 232, 231, 232, 233, 233, 232, 232, 232, 233, 234, 233, 232, 233, 232, 234, 234, 233, 233, 233, 235, 236, 235, 233, 234, 235, 237, 236, 235, 231, 221, 166, 108, 102, 96, 98, 90, 91, 91, 90, 92, 118, 98, 82, 85, 82, 83, 75, 83, 80, 83, 80, 96, 86, 85, 81, 78, 79, 75, 79, 80, 85, 76, 81, 103, 100, 83, 81, 77, 75, 81, 78, 80, 75, 77, 81, 85, 98, 91, 85, 77, 76, 72, 81, 75, 74, 73, 69, 74, 68, 93, 84, 74, 73, 65, 68, 69, 65, 64, 70, 70, 64, 69, 76, 84, 104, 109, 104, 116, 103, 94, 83, 62, 60, 64, 70, 65, 73, 74, 79, 92, 95, 101, 112, 110, 115, 115, 109, 110, 104, 106, 103, 100, 105, 108, 106, 102, 104, 104, 95, 100, 100, 103, 103, 105, 105, 104, 99, 102, 204, 200, 203, 206, 140, 202, 210, 211, 210, 204, 204, 200, 188, 108, 94, 101, 95, 97, 98, 97, 94, 97, 95, 105, 149, 88, 88, 112, 165, 160, 111, 97, 94, 96, 97, 91, 94, 112, 136, 156, 139, 154, 171, 175, 167, 155, 126, 99, 128, 149, 169, 161, 166, 191, 161, 184, 184, 149, 156, 131, 127, 128, 131, 135, 135, 146, 137, 138, 139, 141, 137, 143, 139, 141, 145, 138, 138, 143, 146, 145, 148, 156, 160, 168, 191, 193, 215, 188, 126, 158, 124, 152, 227, 231, 231, 231, 232, 231, 230, 231, 232, 232, 231, 231, 231, 232, 233, 233, 232, 232, 231, 233, 233, 232, 232, 232, 233, 234, 233, 233, 232, 231, 234, 234, 233, 234, 234, 236, 236, 235, 233, 234, 233, 236, 236, 232, 231, 221, 157, 103, 106, 95, 94, 92, 91, 92, 89, 93, 115, 95, 91, 86, 78, 81, 86, 84, 80, 81, 77, 99, 89, 83, 84, 82, 82, 79, 82, 79, 81, 76, 88, 99, 97, 82, 76, 82, 80, 82, 80, 76, 81, 74, 80, 94, 97, 93, 84, 79, 78, 78, 79, 75, 78, 71, 75, 76, 80, 99, 90, 82, 70, 76, 65, 72, 68, 62, 69, 72, 69, 74, 75, 80, 89, 99, 112, 103, 94, 91, 79, 79, 73, 79, 97, 101, 105, 102, 111, 106, 102, 109, 107, 107, 107, 109, 109, 101, 103, 106, 111, 107, 105, 102, 103, 107, 109, 101, 98, 100, 99, 98, 98, 100, 102, 101, 98, 100, 202, 203, 202, 205, 129, 205, 208, 209, 205, 206, 204, 196, 191, 112, 94, 96, 97, 94, 100, 92, 92, 96, 96, 101, 142, 88, 94, 132, 164, 160, 116, 103, 102, 101, 96, 97, 103, 103, 144, 153, 147, 173, 181, 179, 176, 158, 139, 100, 131, 154, 170, 153, 161, 187, 165, 179, 179, 151, 146, 134, 141, 143, 148, 150, 155, 149, 141, 140, 147, 143, 139, 145, 140, 144, 143, 142, 139, 140, 139, 146, 153, 153, 158, 171, 189, 191, 208, 176, 130, 159, 124, 153, 226, 230, 230, 232, 231, 230, 230, 231, 231, 232, 231, 231, 231, 232, 232, 232, 232, 232, 232, 233, 233, 232, 232, 232, 233, 234, 233, 232, 232, 232, 234, 233, 233, 234, 234, 234, 235, 233, 231, 234, 234, 237, 237, 231, 231, 219, 149, 109, 103, 97, 98, 101, 96, 90, 93, 97, 108, 96, 89, 84, 81, 84, 86, 85, 85, 80, 81, 96, 82, 84, 85, 84, 90, 85, 82, 82, 90, 83, 92, 98, 98, 89, 80, 80, 83, 83, 81, 80, 77, 77, 86, 99, 104, 94, 90, 97, 78, 79, 83, 76, 80, 82, 87, 85, 82, 93, 87, 87, 78, 76, 69, 77, 69, 75, 73, 72, 74, 67, 84, 72, 90, 84, 95, 93, 109, 110, 103, 98, 102, 107, 107, 107, 101, 107, 105, 100, 104, 102, 99, 100, 102, 109, 105, 103, 98, 99, 106, 105, 105, 103, 102, 103, 107, 107, 106, 101, 107, 103, 103, 97, 101, 108, 103, 103, 201, 202, 200, 204, 138, 206, 212, 210, 205, 205, 208, 200, 191, 106, 97, 94, 94, 98, 102, 97, 96, 98, 96, 102, 137, 94, 95, 135, 153, 153, 111, 106, 109, 107, 100, 100, 100, 110, 162, 160, 151, 174, 183, 180, 175, 162, 139, 103, 129, 150, 163, 152, 156, 188, 161, 182, 176, 155, 153, 147, 149, 155, 157, 163, 161, 150, 144, 145, 147, 143, 142, 146, 144, 146, 146, 145, 145, 145, 142, 154, 158, 164, 165, 176, 190, 194, 199, 158, 125, 155, 126, 154, 227, 230, 231, 231, 231, 230, 230, 230, 232, 232, 231, 231, 231, 232, 232, 232, 232, 232, 232, 233, 233, 233, 232, 231, 233, 234, 233, 232, 230, 232, 234, 231, 233, 232, 233, 232, 235, 231, 231, 231, 232, 232, 236, 229, 227, 218, 148, 116, 113, 114, 104, 109, 104, 101, 101, 103, 116, 103, 88, 88, 83, 82, 83, 84, 79, 87, 85, 99, 94, 86, 86, 87, 89, 91, 84, 89, 86, 86, 90, 102, 95, 87, 81, 83, 84, 85, 82, 82, 90, 85, 88, 105, 107, 95, 100, 93, 92, 87, 84, 81, 83, 79, 96, 99, 94, 112, 91, 94, 83, 81, 78, 79, 79, 78, 81, 75, 81, 80, 80, 78, 98, 89, 88, 90, 107, 114, 109, 105, 114, 106, 106, 105, 107, 104, 101, 110, 102, 109, 99, 105, 102, 102, 107, 102, 99, 102, 104, 106, 101, 104, 104, 99, 105, 103, 101, 99, 106, 106, 96, 101, 101, 102, 100, 105, 199, 204, 203, 204, 146, 203, 210, 208, 208, 203, 203, 197, 186, 113, 96, 94, 94, 95, 104, 99, 97, 99, 93, 103, 127, 94, 83, 93, 103, 109, 115, 109, 109, 115, 111, 102, 109, 134, 168, 164, 164, 172, 177, 182, 172, 167, 137, 100, 130, 156, 162, 149, 160, 184, 164, 184, 184, 155, 156, 155, 165, 165, 167, 171, 169, 151, 144, 148, 150, 146, 148, 142, 147, 144, 140, 152, 152, 162, 155, 158, 156, 157, 167, 176, 192, 195, 191, 154, 129, 157, 125, 152, 227, 230, 231, 231, 231, 231, 230, 231, 232, 232, 232, 231, 231, 232, 233, 233, 232, 231, 232, 233, 233, 233, 232, 231, 232, 231, 232, 232, 227, 229, 231, 230, 231, 231, 231, 232, 234, 232, 232, 229, 228, 231, 234, 231, 225, 219, 151, 113, 113, 114, 107, 109, 110, 101, 106, 105, 116, 102, 99, 91, 91, 90, 88, 92, 85, 88, 90, 97, 96, 99, 86, 89, 90, 92, 85, 88, 86, 92, 92, 106, 102, 95, 81, 82, 89, 84, 86, 84, 87, 85, 96, 103, 99, 108, 97, 98, 92, 90, 91, 84, 91, 85, 105, 106, 92, 109, 89, 95, 87, 89, 80, 84, 83, 85, 89, 91, 84, 83, 83, 86, 115, 97, 97, 100, 113, 118, 111, 109, 106, 109, 106, 111, 108, 115, 109, 106, 105, 113, 102, 111, 106, 113, 114, 110, 106, 106, 105, 104, 109, 105, 99, 101, 103, 103, 96, 99, 99, 98, 94, 101, 102, 96, 101, 99, 197, 201, 199, 203, 132, 198, 206, 207, 208, 204, 200, 196, 182, 104, 104, 100, 91, 102, 107, 103, 99, 104, 106, 104, 124, 87, 84, 77, 87, 81, 126, 122, 115, 107, 105, 96, 105, 141, 164, 161, 159, 170, 180, 180, 171, 167, 137, 102, 131, 153, 159, 140, 162, 179, 171, 185, 182, 159, 152, 159, 169, 164, 165, 167, 163, 148, 144, 144, 141, 140, 140, 142, 136, 140, 139, 144, 153, 161, 159, 166, 164, 167, 168, 175, 194, 190, 177, 149, 139, 155, 132, 160, 228, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 233, 232, 232, 231, 232, 233, 233, 232, 231, 231, 232, 231, 232, 231, 226, 229, 231, 230, 229, 232, 230, 231, 231, 233, 232, 228, 227, 232, 233, 228, 227, 216, 150, 117, 119, 122, 113, 115, 115, 109, 110, 110, 116, 107, 98, 92, 98, 86, 93, 95, 94, 97, 92, 103, 100, 94, 96, 86, 90, 93, 87, 85, 87, 84, 97, 99, 104, 98, 87, 88, 93, 86, 90, 89, 90, 95, 94, 105, 96, 105, 100, 103, 95, 100, 93, 89, 97, 97, 98, 104, 89, 112, 96, 99, 89, 85, 86, 82, 87, 87, 85, 87, 85, 83, 87, 95, 108, 109, 94, 100, 113, 117, 114, 108, 108, 104, 108, 107, 110, 117, 110, 115, 108, 107, 108, 104, 109, 109, 111, 104, 102, 106, 100, 101, 107, 104, 110, 103, 100, 107, 101, 103, 93, 101, 99, 101, 97, 94, 94, 95, 198, 199, 197, 200, 144, 195, 208, 206, 210, 208, 197, 197, 180, 107, 104, 102, 93, 109, 108, 96, 101, 99, 100, 110, 125, 95, 83, 80, 90, 85, 119, 137, 124, 111, 106, 112, 124, 142, 175, 157, 162, 168, 174, 178, 171, 165, 139, 106, 138, 145, 153, 136, 164, 181, 178, 183, 182, 166, 152, 145, 148, 143, 144, 140, 137, 134, 130, 129, 131, 129, 122, 131, 122, 128, 140, 144, 147, 152, 161, 163, 163, 167, 169, 178, 191, 193, 171, 148, 139, 161, 133, 158, 228, 230, 232, 232, 231, 231, 231, 231, 232, 232, 231, 231, 230, 232, 232, 232, 232, 231, 231, 232, 233, 233, 231, 231, 231, 232, 232, 231, 228, 230, 232, 229, 226, 231, 230, 231, 233, 232, 229, 230, 227, 231, 234, 229, 223, 215, 144, 124, 142, 125, 124, 120, 119, 113, 112, 112, 117, 107, 100, 103, 100, 95, 92, 95, 98, 103, 96, 104, 101, 89, 96, 91, 93, 90, 86, 91, 96, 86, 104, 103, 105, 94, 95, 86, 91, 89, 91, 89, 86, 92, 97, 112, 100, 110, 109, 95, 94, 99, 104, 101, 97, 97, 107, 102, 102, 109, 102, 97, 91, 92, 86, 84, 88, 93, 91, 93, 82, 87, 88, 97, 110, 113, 89, 102, 111, 109, 108, 102, 108, 101, 109, 112, 112, 114, 110, 113, 114, 111, 104, 105, 103, 110, 113, 107, 106, 103, 103, 103, 110, 105, 106, 107, 102, 101, 102, 102, 104, 105, 103, 103, 105, 98, 107, 106, 201, 196, 197, 203, 127, 200, 207, 208, 205, 208, 203, 191, 175, 107, 102, 108, 99, 115, 110, 100, 101, 102, 104, 115, 125, 96, 85, 85, 86, 88, 116, 134, 137, 125, 120, 126, 138, 156, 155, 151, 156, 159, 176, 175, 169, 168, 145, 106, 128, 144, 166, 141, 156, 184, 172, 178, 179, 178, 161, 150, 144, 138, 138, 137, 133, 130, 126, 124, 126, 123, 126, 123, 131, 133, 136, 142, 148, 156, 160, 162, 170, 167, 172, 180, 191, 189, 169, 155, 141, 156, 135, 166, 228, 230, 232, 232, 231, 230, 230, 230, 232, 232, 231, 231, 230, 232, 232, 232, 231, 231, 232, 232, 233, 232, 231, 231, 231, 231, 231, 230, 228, 229, 230, 228, 228, 230, 229, 231, 230, 230, 228, 228, 227, 229, 229, 227, 220, 216, 144, 127, 144, 125, 121, 119, 118, 117, 115, 115, 119, 114, 107, 103, 100, 101, 97, 101, 99, 104, 103, 105, 102, 97, 95, 93, 89, 93, 94, 96, 89, 96, 102, 108, 105, 101, 94, 97, 91, 95, 90, 92, 93, 89, 94, 110, 105, 108, 102, 102, 103, 93, 107, 106, 100, 108, 109, 101, 97, 118, 101, 98, 103, 91, 87, 91, 90, 91, 94, 93, 91, 90, 98, 101, 117, 120, 95, 106, 108, 115, 114, 104, 104, 113, 111, 115, 110, 110, 109, 108, 114, 112, 108, 112, 110, 115, 110, 117, 111, 108, 113, 102, 113, 113, 102, 110, 112, 110, 109, 108, 107, 110, 107, 109, 110, 103, 115, 110, 196, 198, 200, 204, 118, 202, 207, 205, 211, 205, 201, 191, 174, 109, 102, 102, 100, 122, 106, 104, 102, 114, 109, 123, 125, 102, 87, 82, 84, 93, 118, 134, 128, 111, 110, 115, 110, 130, 120, 130, 133, 140, 172, 175, 168, 172, 141, 105, 134, 148, 179, 148, 156, 167, 169, 184, 181, 184, 172, 166, 157, 157, 157, 154, 149, 142, 134, 136, 134, 128, 128, 131, 132, 135, 143, 144, 159, 162, 172, 171, 170, 173, 175, 186, 193, 189, 167, 154, 140, 153, 140, 169, 228, 230, 232, 232, 231, 231, 230, 230, 232, 231, 231, 231, 231, 232, 232, 232, 231, 231, 231, 232, 232, 231, 231, 230, 231, 230, 229, 229, 227, 228, 229, 228, 228, 225, 225, 230, 229, 230, 227, 227, 226, 227, 228, 227, 219, 214, 150, 126, 131, 128, 127, 121, 120, 121, 120, 118, 120, 116, 114, 112, 105, 103, 102, 104, 105, 107, 106, 112, 105, 100, 94, 93, 98, 93, 96, 94, 100, 95, 100, 110, 104, 98, 98, 99, 99, 97, 95, 98, 94, 97, 108, 118, 104, 108, 113, 99, 103, 97, 94, 94, 100, 110, 103, 107, 99, 113, 101, 100, 90, 90, 87, 90, 91, 89, 95, 94, 92, 92, 96, 112, 122, 124, 101, 110, 120, 123, 119, 107, 104, 110, 102, 113, 114, 116, 115, 117, 118, 117, 123, 122, 120, 117, 124, 117, 116, 119, 112, 108, 116, 116, 110, 112, 111, 112, 106, 111, 104, 108, 111, 110, 111, 105, 113, 112, 202, 202, 200, 203, 139, 205, 208, 205, 207, 203, 203, 196, 176, 111, 100, 106, 98, 116, 112, 110, 107, 111, 114, 120, 125, 114, 92, 85, 89, 89, 117, 135, 121, 106, 109, 106, 101, 108, 116, 132, 136, 128, 166, 167, 172, 169, 138, 112, 133, 154, 177, 138, 161, 155, 173, 190, 187, 190, 187, 177, 179, 169, 171, 171, 161, 159, 147, 149, 141, 135, 134, 137, 151, 148, 140, 155, 160, 171, 176, 176, 178, 181, 179, 192, 191, 189, 172, 144, 141, 157, 139, 168, 228, 230, 232, 232, 231, 230, 230, 231, 232, 231, 231, 231, 231, 232, 232, 232, 231, 231, 231, 232, 232, 231, 230, 228, 229, 227, 230, 228, 228, 228, 230, 228, 228, 227, 224, 226, 229, 231, 228, 228, 226, 226, 227, 223, 219, 213, 151, 130, 126, 131, 127, 124, 130, 125, 115, 128, 127, 118, 115, 110, 107, 100, 102, 103, 110, 106, 107, 117, 108, 100, 99, 98, 101, 103, 93, 92, 96, 96, 100, 105, 107, 102, 97, 98, 95, 100, 97, 97, 98, 97, 100, 120, 107, 111, 111, 108, 107, 97, 117, 104, 102, 104, 116, 102, 100, 126, 105, 104, 96, 95, 96, 95, 96, 98, 95, 92, 98, 95, 101, 113, 124, 125, 98, 115, 118, 118, 115, 107, 111, 111, 117, 112, 119, 114, 118, 112, 118, 118, 127, 120, 120, 116, 120, 117, 120, 119, 112, 110, 114, 109, 113, 119, 114, 113, 115, 105, 107, 108, 112, 105, 110, 113, 111, 114, 200, 201, 201, 199, 128, 204, 205, 203, 204, 199, 202, 196, 165, 110, 94, 108, 104, 113, 112, 117, 114, 114, 123, 119, 129, 117, 96, 88, 91, 91, 120, 131, 111, 114, 118, 108, 102, 105, 111, 129, 130, 124, 140, 165, 166, 165, 138, 116, 140, 148, 178, 138, 151, 151, 174, 191, 189, 191, 189, 188, 189, 183, 184, 183, 174, 172, 164, 160, 154, 139, 137, 138, 159, 162, 170, 180, 177, 182, 189, 191, 193, 196, 196, 202, 192, 190, 167, 147, 137, 152, 135, 163, 227, 230, 231, 232, 232, 230, 230, 231, 232, 232, 232, 231, 231, 232, 232, 231, 231, 231, 230, 231, 232, 228, 230, 227, 228, 228, 230, 228, 227, 229, 228, 227, 227, 225, 225, 228, 228, 230, 223, 226, 226, 220, 226, 223, 219, 213, 146, 134, 132, 131, 133, 123, 125, 123, 121, 124, 128, 119, 115, 114, 113, 106, 106, 105, 105, 105, 103, 113, 113, 105, 105, 99, 101, 105, 101, 95, 99, 105, 104, 110, 109, 105, 106, 98, 101, 107, 101, 102, 103, 105, 103, 120, 110, 111, 117, 100, 103, 100, 119, 104, 108, 106, 116, 107, 103, 123, 107, 103, 101, 98, 103, 97, 94, 100, 99, 102, 91, 96, 104, 116, 124, 115, 103, 116, 118, 121, 122, 115, 114, 112, 115, 116, 115, 111, 114, 112, 118, 117, 113, 116, 116, 118, 124, 121, 114, 116, 115, 110, 114, 109, 112, 110, 114, 116, 116, 111, 107, 113, 112, 110, 111, 111, 115, 109, 198, 198, 196, 203, 126, 200, 202, 204, 201, 202, 198, 197, 159, 114, 106, 112, 110, 122, 115, 121, 113, 111, 118, 122, 133, 129, 108, 97, 98, 103, 120, 131, 130, 130, 132, 117, 113, 109, 119, 129, 139, 118, 123, 147, 157, 161, 138, 121, 135, 150, 176, 134, 151, 148, 174, 188, 185, 189, 191, 190, 187, 187, 190, 188, 187, 181, 177, 165, 157, 147, 144, 140, 160, 172, 183, 190, 196, 196, 198, 204, 201, 204, 203, 206, 198, 192, 163, 150, 142, 147, 136, 162, 226, 230, 231, 232, 231, 230, 230, 231, 232, 231, 232, 230, 231, 231, 231, 231, 230, 231, 231, 231, 229, 226, 228, 229, 228, 228, 230, 227, 225, 225, 226, 228, 225, 223, 225, 224, 224, 228, 225, 227, 225, 224, 225, 224, 219, 213, 148, 138, 132, 130, 127, 130, 129, 126, 126, 130, 125, 122, 114, 114, 115, 112, 110, 110, 116, 110, 107, 115, 113, 112, 109, 106, 108, 106, 106, 103, 99, 105, 105, 111, 108, 111, 109, 104, 108, 103, 103, 107, 105, 106, 103, 122, 105, 114, 114, 109, 111, 108, 118, 110, 116, 111, 118, 117, 105, 130, 112, 108, 105, 101, 105, 102, 98, 100, 99, 99, 98, 101, 108, 121, 121, 125, 103, 112, 122, 116, 111, 116, 112, 116, 115, 117, 112, 120, 122, 118, 120, 121, 124, 120, 125, 126, 124, 120, 122, 115, 115, 115, 119, 117, 115, 106, 115, 111, 113, 111, 109, 120, 113, 111, 116, 112, 113, 113, 197, 193, 193, 199, 124, 199, 202, 201, 202, 198, 199, 192, 155, 108, 105, 109, 117, 131, 116, 115, 122, 117, 124, 135, 145, 141, 112, 102, 102, 112, 121, 142, 158, 156, 154, 129, 128, 123, 123, 121, 122, 121, 120, 124, 154, 158, 140, 121, 135, 148, 168, 142, 149, 148, 173, 186, 189, 189, 189, 191, 190, 190, 194, 192, 189, 190, 187, 176, 160, 152, 146, 145, 152, 179, 192, 194, 196, 203, 198, 209, 207, 207, 205, 206, 197, 189, 161, 154, 143, 153, 133, 161, 224, 230, 231, 230, 230, 229, 230, 230, 231, 231, 231, 231, 231, 231, 232, 232, 231, 231, 231, 231, 231, 226, 228, 225, 228, 228, 230, 226, 226, 226, 227, 228, 226, 223, 224, 224, 225, 225, 225, 225, 223, 225, 225, 223, 220, 217, 152, 138, 134, 129, 129, 126, 131, 126, 125, 126, 131, 122, 114, 114, 112, 106, 111, 112, 113, 112, 107, 118, 115, 110, 109, 108, 110, 104, 104, 114, 105, 109, 107, 113, 115, 112, 107, 104, 110, 109, 107, 112, 107, 106, 106, 127, 116, 115, 117, 115, 115, 111, 115, 107, 115, 107, 122, 112, 106, 132, 110, 113, 103, 102, 102, 107, 101, 104, 112, 106, 102, 101, 106, 123, 120, 119, 103, 119, 113, 118, 120, 120, 112, 120, 123, 121, 117, 121, 118, 122, 124, 123, 124, 118, 120, 122, 123, 116, 125, 119, 112, 118, 116, 115, 118, 111, 113, 114, 115, 112, 108, 109, 111, 118, 115, 114, 114, 115, 198, 192, 191, 194, 135, 198, 198, 198, 202, 197, 195, 190, 151, 111, 109, 117, 122, 137, 122, 120, 134, 124, 131, 133, 156, 146, 105, 101, 104, 124, 125, 152, 165, 165, 158, 135, 127, 125, 128, 118, 109, 113, 113, 123, 139, 158, 141, 111, 132, 150, 153, 136, 149, 144, 175, 192, 192, 195, 193, 190, 191, 194, 195, 192, 193, 193, 192, 185, 176, 152, 150, 150, 149, 180, 191, 192, 198, 201, 201, 206, 204, 205, 204, 203, 191, 190, 164, 161, 142, 156, 144, 162, 223, 230, 231, 231, 231, 230, 230, 231, 232, 230, 230, 230, 231, 232, 231, 230, 230, 230, 230, 231, 230, 229, 228, 224, 227, 230, 230, 227, 227, 227, 229, 224, 224, 224, 222, 225, 224, 225, 225, 226, 226, 224, 223, 223, 221, 212, 162, 137, 135, 129, 133, 127, 132, 129, 126, 126, 129, 125, 125, 113, 115, 110, 109, 117, 112, 105, 109, 120, 113, 114, 113, 106, 108, 113, 106, 102, 105, 108, 106, 116, 115, 110, 106, 108, 112, 109, 111, 103, 105, 108, 106, 124, 112, 117, 115, 115, 117, 117, 115, 114, 114, 115, 121, 117, 112, 134, 117, 117, 110, 119, 115, 101, 104, 107, 110, 105, 125, 109, 111, 125, 120, 123, 108, 122, 117, 118, 123, 115, 121, 118, 117, 123, 123, 114, 125, 125, 125, 124, 121, 122, 125, 126, 122, 123, 124, 120, 117, 120, 113, 114, 122, 108, 114, 114, 112, 115, 111, 111, 112, 117, 117, 113, 115, 111, 193, 193, 189, 199, 130, 195, 196, 195, 201, 196, 198, 189, 148, 114, 114, 121, 122, 156, 152, 147, 145, 132, 133, 140, 174, 156, 107, 106, 115, 125, 122, 157, 164, 159, 153, 144, 128, 129, 128, 123, 109, 111, 111, 122, 128, 150, 137, 113, 128, 155, 155, 135, 157, 147, 179, 187, 191, 193, 193, 192, 198, 195, 197, 197, 199, 193, 192, 182, 176, 154, 150, 146, 159, 168, 192, 192, 197, 201, 203, 205, 208, 206, 205, 200, 192, 192, 162, 161, 143, 155, 138, 163, 218, 230, 231, 231, 231, 230, 230, 230, 231, 231, 229, 228, 230, 231, 231, 231, 227, 228, 228, 229, 228, 229, 224, 226, 224, 227, 228, 222, 228, 224, 228, 226, 225, 223, 223, 222, 222, 224, 224, 222, 222, 222, 222, 220, 220, 208, 162, 143, 139, 141, 130, 132, 132, 130, 131, 131, 132, 128, 117, 117, 117, 116, 115, 112, 112, 107, 112, 119, 118, 114, 115, 117, 108, 109, 108, 108, 113, 111, 105, 123, 122, 107, 107, 109, 109, 113, 105, 106, 106, 108, 108, 130, 120, 117, 116, 114, 116, 116, 132, 122, 117, 118, 128, 123, 121, 129, 118, 122, 112, 118, 111, 110, 109, 112, 112, 107, 103, 107, 110, 124, 125, 131, 112, 116, 118, 126, 124, 119, 122, 120, 118, 115, 122, 121, 117, 123, 121, 124, 124, 123, 122, 126, 122, 131, 125, 124, 119, 124, 117, 116, 117, 116, 122, 120, 113, 115, 119, 112, 124, 115, 115, 116, 116, 114, 197, 191, 191, 193, 112, 186, 194, 199, 193, 195, 194, 188, 148, 111, 112, 121, 129, 165, 162, 160, 153, 132, 136, 149, 168, 162, 113, 109, 129, 128, 114, 148, 165, 160, 152, 141, 134, 134, 137, 131, 115, 108, 113, 110, 113, 135, 137, 115, 136, 157, 155, 140, 160, 149, 178, 193, 193, 191, 189, 196, 193, 196, 193, 198, 197, 194, 194, 189, 180, 165, 156, 150, 158, 166, 187, 192, 193, 198, 198, 204, 206, 206, 206, 196, 194, 195, 165, 168, 146, 153, 144, 166, 223, 228, 229, 230, 231, 229, 229, 230, 227, 231, 230, 230, 229, 229, 231, 231, 226, 227, 228, 230, 231, 228, 222, 226, 223, 223, 224, 225, 224, 222, 224, 225, 225, 222, 222, 223, 221, 224, 226, 221, 221, 225, 216, 224, 219, 210, 166, 141, 140, 134, 132, 135, 132, 130, 133, 130, 135, 125, 127, 122, 118, 113, 118, 116, 116, 117, 117, 124, 119, 120, 120, 123, 121, 111, 118, 120, 117, 117, 115, 116, 118, 113, 112, 109, 110, 112, 114, 113, 109, 108, 108, 129, 120, 121, 124, 123, 126, 124, 133, 124, 124, 118, 124, 126, 128, 134, 120, 118, 118, 110, 116, 110, 113, 110, 112, 111, 108, 112, 109, 126, 122, 133, 115, 117, 122, 124, 122, 123, 121, 124, 121, 121, 125, 120, 118, 126, 127, 132, 125, 122, 128, 125, 131, 126, 124, 128, 122, 129, 117, 119, 121, 124, 121, 130, 124, 127, 117, 122, 125, 122, 128, 126, 122, 115, 192, 190, 194, 192, 113, 186, 195, 193, 194, 194, 197, 184, 146, 122, 112, 128, 132, 162, 167, 164, 157, 138, 145, 163, 182, 169, 121, 129, 127, 127, 116, 146, 148, 155, 142, 137, 132, 128, 140, 138, 121, 115, 110, 117, 122, 130, 138, 120, 143, 157, 155, 141, 155, 149, 177, 190, 196, 195, 189, 193, 195, 190, 193, 199, 196, 195, 192, 190, 177, 169, 158, 159, 157, 163, 187, 194, 197, 197, 202, 202, 202, 202, 198, 192, 192, 186, 171, 166, 144, 152, 152, 165, 222, 228, 231, 230, 231, 229, 229, 229, 230, 230, 229, 230, 229, 229, 230, 228, 226, 229, 227, 228, 230, 226, 222, 223, 224, 226, 226, 227, 224, 225, 224, 226, 225, 225, 220, 222, 224, 226, 225, 226, 221, 224, 222, 220, 219, 210, 172, 148, 142, 145, 140, 133, 137, 135, 138, 131, 133, 135, 129, 129, 118, 115, 116, 120, 122, 116, 120, 122, 122, 125, 117, 115, 118, 116, 123, 122, 120, 115, 116, 125, 123, 120, 112, 117, 119, 115, 117, 117, 116, 119, 115, 126, 131, 128, 124, 120, 125, 119, 122, 124, 126, 118, 128, 124, 121, 137, 127, 121, 114, 112, 114, 112, 112, 112, 117, 107, 107, 114, 113, 124, 131, 134, 123, 124, 127, 128, 134, 129, 126, 122, 123, 125, 128, 127, 122, 125, 129, 130, 127, 126, 132, 128, 130, 128, 125, 131, 126, 132, 126, 123, 128, 130, 130, 127, 126, 125, 122, 123, 128, 123, 122, 123, 116, 120, 194, 187, 190, 196, 109, 187, 191, 195, 191, 191, 193, 186, 142, 123, 111, 124, 132, 161, 168, 170, 162, 162, 167, 178, 183, 172, 145, 132, 126, 133, 121, 137, 138, 140, 131, 124, 118, 116, 137, 128, 121, 124, 116, 121, 122, 123, 143, 124, 143, 161, 153, 142, 152, 148, 178, 193, 194, 192, 197, 193, 193, 199, 192, 199, 198, 193, 195, 189, 177, 170, 156, 156, 157, 166, 178, 190, 197, 197, 200, 202, 203, 203, 200, 193, 192, 188, 167, 156, 142, 162, 147, 168, 219, 227, 231, 231, 231, 230, 230, 229, 229, 230, 229, 228, 229, 230, 230, 226, 226, 225, 219, 225, 229, 227, 226, 222, 224, 224, 224, 224, 222, 223, 223, 221, 223, 222, 220, 223, 222, 221, 224, 222, 219, 219, 221, 217, 219, 211, 184, 149, 147, 143, 146, 143, 145, 145, 140, 138, 140, 135, 142, 134, 128, 128, 121, 127, 122, 124, 124, 126, 132, 128, 122, 123, 117, 122, 129, 123, 121, 116, 122, 125, 126, 126, 121, 118, 119, 123, 122, 119, 119, 124, 123, 127, 132, 133, 127, 127, 128, 122, 134, 121, 121, 119, 125, 129, 127, 142, 124, 128, 116, 118, 116, 117, 129, 117, 115, 117, 112, 111, 121, 124, 135, 129, 119, 128, 128, 129, 135, 131, 127, 134, 125, 129, 128, 126, 127, 132, 130, 129, 132, 127, 126, 132, 129, 129, 128, 131, 135, 131, 130, 127, 123, 129, 130, 126, 126, 125, 126, 123, 125, 122, 121, 124, 116, 118, 193, 187, 189, 193, 116, 191, 192, 193, 195, 194, 184, 184, 145, 119, 110, 127, 143, 167, 169, 169, 169, 173, 172, 180, 181, 177, 146, 131, 126, 136, 123, 132, 133, 134, 124, 116, 120, 119, 132, 135, 123, 130, 123, 123, 125, 124, 140, 126, 147, 158, 154, 142, 155, 151, 177, 190, 196, 192, 194, 192, 192, 199, 198, 200, 197, 194, 191, 188, 170, 168, 158, 157, 159, 164, 173, 190, 192, 198, 199, 202, 201, 200, 198, 190, 188, 184, 165, 155, 150, 159, 155, 168, 224, 229, 231, 231, 230, 229, 230, 228, 228, 229, 228, 230, 229, 228, 228, 227, 225, 225, 228, 225, 228, 227, 226, 221, 224, 224, 223, 223, 225, 223, 223, 223, 223, 222, 221, 220, 222, 222, 222, 216, 220, 216, 216, 221, 216, 210, 185, 158, 154, 151, 151, 150, 150, 152, 150, 142, 150, 141, 147, 140, 132, 132, 123, 127, 129, 127, 122, 126, 128, 129, 127, 124, 119, 118, 125, 126, 128, 121, 119, 131, 132, 129, 132, 123, 124, 121, 129, 127, 137, 135, 125, 130, 138, 130, 120, 130, 125, 131, 138, 134, 126, 126, 137, 133, 129, 149, 134, 131, 121, 121, 123, 123, 124, 120, 116, 119, 114, 118, 119, 130, 134, 130, 121, 129, 128, 131, 133, 131, 128, 131, 132, 135, 135, 131, 136, 128, 134, 134, 133, 133, 135, 136, 134, 133, 130, 133, 136, 132, 128, 128, 131, 132, 128, 129, 128, 127, 122, 126, 120, 125, 126, 125, 126, 122, 186, 188, 188, 192, 111, 188, 192, 197, 193, 192, 190, 182, 139, 111, 111, 128, 144, 169, 168, 171, 166, 172, 177, 182, 187, 183, 147, 120, 133, 120, 115, 121, 125, 126, 121, 119, 114, 119, 127, 135, 118, 127, 122, 131, 122, 125, 144, 129, 143, 155, 150, 145, 154, 154, 178, 192, 195, 196, 190, 194, 194, 196, 195, 195, 197, 196, 198, 191, 179, 173, 160, 157, 158, 161, 167, 178, 195, 196, 199, 198, 198, 202, 192, 190, 191, 176, 160, 155, 148, 160, 155, 170, 221, 228, 228, 228, 229, 228, 229, 230, 229, 229, 228, 229, 229, 228, 229, 226, 226, 227, 229, 226, 227, 228, 225, 224, 224, 224, 224, 223, 226, 220, 226, 223, 221, 220, 219, 220, 221, 221, 221, 223, 222, 219, 216, 221, 216, 214, 195, 162, 163, 162, 157, 156, 156, 153, 155, 157, 150, 147, 149, 143, 130, 131, 128, 128, 133, 129, 128, 126, 126, 131, 131, 130, 123, 120, 131, 127, 132, 135, 131, 135, 128, 128, 130, 128, 135, 132, 128, 123, 136, 130, 132, 127, 135, 136, 126, 133, 134, 136, 134, 137, 131, 128, 136, 142, 130, 142, 137, 137, 129, 130, 131, 134, 131, 127, 126, 118, 121, 124, 125, 132, 141, 142, 128, 130, 138, 140, 137, 134, 135, 138, 136, 133, 137, 137, 133, 135, 138, 135, 138, 130, 134, 137, 133, 131, 135, 141, 136, 134, 135, 134, 130, 136, 124, 130, 127, 129, 124, 127, 125, 121, 122, 128, 129, 124, 190, 190, 188, 193, 116, 193, 195, 194, 189, 188, 189, 179, 135, 113, 122, 122, 146, 165, 163, 170, 168, 172, 180, 184, 185, 186, 149, 130, 134, 114, 120, 116, 125, 118, 119, 117, 125, 119, 130, 135, 124, 125, 127, 126, 129, 126, 144, 133, 141, 166, 159, 146, 156, 155, 184, 189, 197, 191, 194, 189, 192, 193, 192, 197, 196, 195, 194, 194, 183, 171, 165, 159, 160, 164, 168, 168, 196, 199, 196, 199, 199, 197, 191, 190, 190, 179, 159, 157, 151, 160, 155, 177, 218, 226, 229, 228, 227, 227, 226, 228, 229, 229, 226, 226, 228, 230, 229, 227, 226, 225, 227, 228, 227, 224, 222, 222, 223, 222, 227, 225, 224, 224, 224, 228, 223, 219, 220, 220, 223, 222, 221, 220, 221, 218, 216, 221, 218, 208, 202, 173, 170, 168, 165, 161, 158, 155, 152, 154, 152, 149, 153, 146, 140, 138, 131, 137, 133, 127, 132, 129, 132, 127, 128, 131, 125, 124, 132, 128, 125, 135, 134, 135, 129, 134, 134, 131, 133, 130, 128, 126, 130, 128, 128, 135, 136, 136, 128, 134, 132, 139, 143, 130, 134, 136, 140, 149, 140, 147, 143, 139, 136, 135, 147, 144, 131, 130, 125, 131, 129, 127, 135, 130, 140, 142, 135, 136, 136, 133, 137, 137, 132, 135, 134, 136, 134, 138, 133, 140, 141, 140, 138, 144, 144, 141, 140, 138, 137, 141, 141, 129, 132, 131, 129, 133, 134, 132, 134, 133, 130, 135, 129, 135, 122, 134, 127, 131, 189, 190, 187, 186, 119, 186, 191, 190, 189, 191, 185, 179, 133, 120, 119, 128, 144, 162, 169, 168, 171, 173, 186, 185, 192, 187, 144, 135, 122, 115, 119, 121, 122, 119, 125, 127, 127, 124, 135, 130, 126, 132, 131, 127, 132, 133, 142, 136, 147, 169, 167, 148, 160, 159, 187, 191, 196, 194, 196, 191, 197, 198, 199, 199, 199, 193, 192, 196, 186, 176, 166, 157, 162, 164, 168, 170, 193, 198, 195, 197, 197, 187, 182, 189, 189, 179, 157, 160, 153, 158, 156, 169, 218, 224, 226, 228, 228, 227, 224, 225, 227, 228, 227, 226, 227, 229, 227, 227, 224, 223, 224, 225, 226, 224, 222, 223, 224, 225, 224, 221, 221, 223, 220, 224, 217, 217, 221, 221, 223, 221, 222, 215, 215, 218, 221, 216, 215, 208, 196, 176, 183, 184, 183, 169, 171, 166, 161, 156, 159, 154, 155, 147, 148, 139, 138, 138, 135, 134, 136, 135, 137, 133, 134, 128, 126, 129, 133, 133, 134, 135, 130, 136, 137, 135, 129, 137, 133, 135, 139, 137, 136, 134, 139, 139, 142, 140, 140, 142, 145, 136, 145, 133, 134, 140, 146, 147, 137, 144, 143, 143, 139, 136, 133, 131, 126, 134, 132, 129, 129, 129, 132, 133, 144, 139, 132, 134, 140, 136, 140, 133, 139, 136, 139, 136, 137, 141, 139, 145, 144, 141, 139, 147, 145, 146, 140, 137, 142, 139, 143, 137, 139, 135, 138, 139, 133, 134, 135, 130, 133, 133, 131, 131, 129, 132, 128, 128, 188, 187, 186, 187, 95, 183, 191, 191, 190, 191, 191, 183, 131, 125, 121, 126, 145, 163, 165, 169, 170, 175, 181, 185, 187, 181, 163, 138, 122, 119, 121, 121, 123, 128, 124, 128, 139, 128, 139, 137, 134, 125, 135, 134, 138, 136, 143, 133, 145, 171, 167, 151, 162, 154, 186, 193, 190, 194, 192, 192, 194, 192, 193, 193, 194, 196, 191, 190, 181, 176, 170, 166, 164, 168, 169, 172, 195, 197, 197, 195, 196, 185, 181, 180, 186, 172, 161, 159, 153, 162, 156, 169, 218, 225, 228, 228, 227, 225, 225, 226, 227, 225, 226, 226, 226, 229, 226, 226, 221, 223, 224, 225, 225, 221, 220, 221, 223, 224, 224, 222, 222, 220, 221, 223, 219, 219, 217, 218, 222, 221, 218, 217, 217, 219, 216, 214, 214, 209, 200, 195, 203, 207, 196, 190, 193, 184, 182, 173, 168, 164, 164, 156, 155, 146, 143, 140, 143, 139, 138, 142, 136, 141, 146, 135, 134, 138, 139, 142, 139, 136, 137, 138, 136, 141, 129, 129, 128, 137, 139, 142, 144, 142, 140, 142, 143, 143, 145, 143, 151, 151, 149, 142, 140, 140, 140, 148, 137, 143, 144, 143, 137, 139, 129, 134, 128, 133, 132, 134, 130, 134, 131, 141, 145, 136, 134, 141, 141, 144, 136, 139, 138, 135, 139, 137, 143, 142, 140, 143, 143, 143, 146, 140, 141, 144, 137, 136, 143, 140, 140, 142, 144, 141, 142, 144, 136, 144, 143, 138, 136, 136, 143, 131, 135, 132, 130, 133, 189, 186, 185, 183, 91, 177, 195, 192, 191, 190, 186, 179, 133, 123, 114, 121, 142, 153, 159, 163, 166, 173, 182, 183, 186, 181, 174, 134, 122, 119, 124, 125, 122, 125, 129, 135, 130, 130, 136, 138, 135, 136, 138, 136, 135, 131, 144, 138, 145, 169, 164, 153, 162, 158, 182, 190, 194, 195, 194, 189, 194, 194, 195, 199, 198, 197, 191, 193, 178, 175, 176, 163, 170, 174, 170, 177, 196, 198, 196, 195, 189, 184, 171, 171, 172, 168, 161, 158, 155, 163, 152, 174, 213, 224, 226, 227, 226, 227, 228, 226, 226, 224, 225, 224, 227, 227, 229, 228, 224, 223, 222, 224, 222, 220, 217, 217, 221, 221, 222, 223, 221, 220, 219, 219, 218, 218, 211, 214, 219, 220, 216, 215, 214, 218, 219, 213, 215, 215, 212, 209, 207, 203, 201, 201, 204, 201, 197, 198, 193, 192, 184, 175, 170, 164, 160, 151, 141, 146, 143, 145, 146, 144, 144, 145, 139, 141, 139, 144, 142, 136, 138, 139, 140, 147, 139, 134, 135, 140, 137, 137, 137, 140, 138, 143, 147, 145, 140, 144, 153, 151, 146, 147, 145, 144, 148, 153, 143, 144, 142, 148, 135, 138, 137, 136, 139, 135, 140, 132, 134, 134, 134, 135, 144, 144, 139, 140, 147, 138, 143, 140, 142, 142, 144, 143, 147, 147, 143, 143, 143, 142, 146, 141, 142, 148, 138, 145, 149, 143, 143, 146, 147, 140, 140, 141, 141, 144, 144, 142, 136, 139, 144, 141, 135, 138, 135, 135, 186, 182, 181, 183, 91, 178, 184, 188, 189, 192, 182, 177, 141, 128, 124, 132, 142, 159, 142, 147, 153, 164, 179, 184, 183, 179, 172, 130, 123, 119, 126, 127, 129, 133, 130, 131, 134, 128, 137, 137, 138, 144, 139, 136, 131, 133, 144, 140, 145, 171, 169, 160, 169, 157, 181, 188, 188, 193, 190, 194, 192, 194, 191, 198, 194, 188, 193, 193, 184, 176, 176, 174, 171, 176, 173, 192, 196, 195, 193, 192, 188, 177, 166, 168, 169, 166, 163, 160, 157, 167, 156, 176, 215, 214, 223, 226, 226, 226, 227, 226, 227, 224, 222, 226, 227, 228, 226, 225, 224, 223, 223, 222, 223, 218, 216, 220, 220, 222, 221, 220, 219, 219, 220, 221, 218, 214, 213, 215, 215, 217, 214, 217, 217, 219, 217, 215, 215, 216, 211, 209, 211, 204, 205, 201, 206, 204, 202, 202, 200, 202, 199, 198, 195, 185, 182, 174, 159, 148, 145, 144, 146, 143, 146, 143, 146, 142, 143, 147, 145, 141, 141, 145, 140, 146, 137, 135, 137, 139, 142, 143, 141, 146, 143, 138, 147, 141, 144, 144, 154, 156, 147, 152, 151, 146, 150, 153, 148, 146, 147, 149, 143, 141, 141, 142, 139, 140, 144, 142, 139, 139, 139, 138, 143, 141, 144, 140, 142, 146, 149, 146, 141, 151, 149, 152, 145, 147, 143, 148, 145, 148, 143, 145, 148, 145, 147, 138, 148, 136, 148, 143, 146, 141, 140, 143, 142, 141, 140, 142, 141, 138, 139, 144, 136, 141, 136, 134, 184, 187, 183, 188, 97, 174, 185, 186, 186, 189, 184, 173, 141, 127, 120, 134, 139, 148, 140, 142, 145, 154, 175, 182, 185, 181, 172, 128, 125, 126, 130, 127, 134, 131, 133, 133, 133, 135, 136, 142, 136, 140, 138, 138, 136, 138, 145, 141, 148, 171, 158, 160, 164, 158, 182, 188, 189, 195, 193, 188, 197, 193, 191, 197, 194, 193, 197, 193, 186, 178, 177, 177, 170, 180, 180, 195, 192, 192, 193, 189, 182, 180, 166, 166, 172, 169, 164, 160, 158, 163, 165, 178, 213, 217, 221, 226, 227, 222, 224, 226, 226, 225, 225, 223, 225, 226, 223, 223, 223, 222, 222, 222, 224, 221, 218, 220, 220, 220, 220, 221, 218, 220, 220, 221, 219, 220, 214, 217, 214, 215, 217, 216, 215, 219, 216, 217, 211, 215, 212, 212, 214, 207, 207, 203, 202, 204, 201, 205, 203, 203, 202, 203, 195, 193, 192, 184, 172, 163, 156, 155, 144, 151, 150, 151, 149, 147, 147, 149, 144, 145, 143, 143, 145, 144, 138, 141, 144, 147, 146, 151, 143, 146, 147, 149, 152, 151, 145, 150, 160, 154, 154, 152, 154, 148, 151, 147, 148, 146, 150, 152, 149, 145, 145, 141, 142, 148, 143, 143, 140, 144, 145, 144, 145, 142, 142, 145, 147, 151, 150, 148, 149, 151, 151, 152, 147, 152, 148, 152, 149, 149, 155, 147, 148, 149, 152, 146, 150, 145, 146, 144, 152, 148, 147, 149, 147, 149, 147, 143, 143, 141, 147, 147, 143, 145, 144, 140, 186, 184, 183, 192, 97, 180, 185, 187, 189, 187, 187, 170, 140, 130, 123, 128, 140, 149, 145, 147, 142, 150, 169, 180, 179, 176, 170, 143, 129, 134, 129, 131, 135, 129, 131, 133, 129, 131, 143, 140, 141, 143, 146, 136, 140, 138, 144, 143, 153, 169, 160, 157, 158, 161, 180, 187, 190, 190, 194, 193, 196, 195, 195, 194, 197, 195, 192, 192, 188, 182, 178, 180, 172, 177, 183, 191, 193, 198, 195, 187, 181, 174, 169, 171, 172, 168, 166, 163, 163, 165, 163, 178, 210, 221, 218, 223, 225, 225, 225, 226, 227, 228, 225, 226, 225, 224, 224, 223, 222, 220, 223, 219, 220, 222, 219, 221, 220, 222, 220, 221, 218, 218, 219, 220, 220, 219, 216, 217, 218, 217, 215, 216, 216, 216, 217, 214, 213, 214, 211, 214, 209, 209, 205, 208, 200, 205, 206, 206, 204, 203, 200, 201, 198, 198, 189, 179, 170, 165, 162, 154, 155, 156, 154, 159, 159, 149, 159, 151, 154, 150, 147, 144, 150, 149, 147, 145, 144, 147, 151, 148, 145, 147, 147, 147, 149, 148, 143, 153, 148, 146, 150, 150, 148, 146, 148, 151, 151, 148, 151, 148, 150, 143, 144, 144, 140, 150, 147, 144, 145, 147, 143, 150, 151, 146, 147, 147, 146, 151, 156, 152, 146, 144, 152, 153, 148, 155, 152, 152, 152, 154, 150, 151, 153, 152, 157, 155, 153, 150, 154, 151, 154, 151, 150, 154, 151, 155, 153, 146, 149, 148, 147, 146, 148, 155, 152, 146, 186, 181, 184, 184, 93, 173, 186, 187, 188, 188, 184, 175, 143, 134, 128, 130, 142, 149, 150, 151, 144, 151, 165, 172, 174, 173, 170, 141, 127, 136, 137, 134, 135, 136, 134, 135, 139, 140, 150, 145, 147, 144, 144, 141, 137, 144, 148, 142, 146, 167, 163, 156, 165, 165, 182, 185, 193, 195, 194, 197, 194, 194, 196, 194, 196, 198, 192, 199, 184, 182, 170, 170, 168, 172, 175, 183, 190, 193, 186, 181, 177, 171, 166, 166, 175, 168, 168, 164, 160, 175, 165, 183, 208, 220, 219, 225, 223, 226, 227, 225, 227, 229, 227, 226, 223, 225, 224, 223, 223, 222, 220, 218, 222, 219, 220, 220, 224, 222, 221, 224, 218, 217, 217, 219, 218, 218, 218, 218, 219, 219, 216, 217, 221, 218, 220, 215, 213, 214, 212, 214, 209, 212, 208, 208, 208, 207, 209, 204, 211, 202, 203, 200, 196, 193, 180, 168, 170, 164, 161, 161, 161, 162, 163, 163, 167, 152, 156, 156, 155, 149, 153, 149, 153, 152, 149, 148, 149, 155, 156, 153, 154, 149, 147, 150, 150, 153, 149, 157, 154, 152, 153, 149, 152, 149, 151, 152, 150, 143, 152, 149, 151, 147, 151, 147, 147, 150, 149, 151, 150, 147, 149, 152, 149, 148, 153, 146, 153, 154, 156, 147, 153, 155, 151, 152, 154, 149, 149, 153, 155, 158, 156, 154, 155, 153, 155, 153, 151, 154, 151, 155, 153, 154, 154, 155, 154, 158, 157, 154, 154, 154, 150, 151, 150, 156, 152, 147, 186, 185, 182, 185, 87, 180, 190, 190, 190, 187, 181, 177, 139, 131, 128, 131, 140, 145, 142, 147, 142, 149, 148, 168, 171, 168, 167, 149, 131, 132, 136, 132, 137, 142, 138, 142, 145, 142, 154, 150, 152, 150, 145, 145, 143, 144, 152, 147, 153, 171, 163, 161, 169, 169, 185, 190, 196, 195, 194, 196, 195, 198, 197, 195, 196, 202, 195, 196, 188, 179, 169, 161, 165, 167, 170, 177, 184, 184, 181, 180, 173, 171, 166, 169, 172, 167, 164, 165, 166, 175, 166, 181, 211, 221, 221, 225, 224, 223, 225, 225, 226, 226, 226, 227, 222, 225, 224, 222, 220, 222, 221, 220, 223, 221, 219, 219, 221, 221, 221, 220, 219, 219, 219, 221, 217, 218, 214, 219, 219, 221, 215, 219, 217, 217, 221, 218, 214, 216, 216, 214, 212, 210, 209, 207, 206, 212, 210, 208, 209, 200, 198, 198, 192, 180, 176, 169, 170, 162, 161, 159, 162, 167, 164, 169, 163, 159, 156, 162, 152, 156, 156, 155, 162, 158, 156, 157, 148, 156, 155, 158, 152, 151, 156, 155, 151, 161, 156, 154, 153, 156, 155, 152, 146, 149, 145, 157, 157, 149, 153, 152, 158, 150, 151, 148, 153, 152, 152, 151, 150, 149, 149, 151, 155, 151, 156, 143, 155, 155, 153, 153, 152, 158, 153, 151, 155, 150, 154, 154, 149, 154, 155, 159, 157, 163, 158, 157, 156, 157, 158, 155, 156, 152, 154, 155, 159, 161, 159, 157, 158, 157, 155, 155, 162, 168, 161, 156, 188, 182, 184, 187, 88, 178, 192, 189, 190, 192, 181, 170, 142, 130, 132, 130, 130, 140, 137, 139, 144, 138, 148, 157, 161, 159, 154, 147, 141, 138, 139, 138, 136, 136, 140, 145, 144, 143, 151, 149, 154, 149, 148, 150, 146, 147, 152, 149, 157, 173, 168, 166, 171, 174, 186, 192, 195, 192, 192, 193, 197, 199, 196, 200, 196, 204, 197, 195, 186, 171, 168, 165, 171, 166, 166, 173, 177, 180, 177, 181, 174, 173, 170, 173, 170, 172, 173, 169, 170, 170, 168, 181, 213, 224, 222, 224, 225, 225, 222, 224, 226, 223, 228, 224, 225, 225, 222, 222, 220, 218, 223, 223, 223, 221, 220, 222, 222, 223, 224, 221, 218, 220, 221, 221, 218, 219, 218, 218, 222, 220, 219, 219, 218, 216, 216, 217, 216, 215, 214, 214, 208, 208, 213, 208, 210, 213, 210, 205, 205, 201, 197, 190, 185, 177, 178, 172, 170, 167, 167, 165, 168, 171, 170, 173, 168, 167, 161, 165, 160, 162, 159, 165, 162, 165, 158, 155, 151, 156, 160, 154, 153, 153, 157, 159, 158, 157, 156, 160, 153, 163, 153, 157, 152, 153, 151, 155, 157, 153, 155, 158, 155, 154, 151, 152, 149, 153, 151, 153, 154, 156, 151, 152, 153, 157, 154, 150, 149, 159, 159, 156, 156, 158, 158, 159, 156, 157, 153, 156, 158, 161, 158, 160, 162, 163, 162, 165, 161, 159, 165, 164, 162, 160, 158, 163, 158, 159, 160, 161, 157, 166, 155, 163, 165, 168, 163, 161, 184, 185, 182, 184, 87, 182, 190, 187, 191, 190, 181, 170, 142, 133, 132, 130, 134, 138, 140, 140, 137, 138, 150, 151, 154, 153, 144, 145, 140, 136, 136, 142, 134, 137, 137, 142, 147, 147, 149, 157, 149, 147, 147, 146, 153, 151, 151, 157, 156, 173, 170, 164, 172, 175, 190, 195, 199, 193, 194, 192, 198, 196, 195, 198, 196, 199, 195, 197, 190, 177, 171, 169, 171, 171, 170, 170, 172, 176, 181, 176, 173, 174, 174, 176, 173, 174, 171, 169, 173, 178, 169, 186, 214, 221, 222, 226, 221, 223, 225, 225, 225, 226, 226, 225, 224, 224, 224, 221, 220, 220, 220, 221, 222, 219, 222, 221, 222, 223, 224, 219, 219, 219, 220, 218, 220, 218, 216, 220, 221, 218, 219, 218, 219, 217, 216, 219, 217, 215, 215, 211, 214, 211, 211, 208, 210, 211, 211, 209, 207, 203, 198, 188, 178, 177, 172, 169, 172, 171, 172, 170, 174, 178, 179, 171, 175, 169, 170, 164, 164, 163, 163, 160, 163, 161, 163, 161, 159, 163, 163, 158, 163, 156, 159, 161, 160, 157, 157, 157, 159, 154, 159, 155, 155, 158, 163, 156, 158, 157, 157, 160, 156, 158, 155, 156, 157, 154, 156, 154, 158, 152, 154, 152, 158, 156, 151, 156, 154, 155, 157, 157, 160, 160, 160, 159, 160, 158, 162, 154, 162, 162, 162, 162, 167, 167, 162, 169, 166, 161, 167, 168, 165, 164, 160, 159, 162, 161, 161, 159, 164, 160, 161, 164, 165, 166, 159, 157, 189, 182, 179, 181, 80, 181, 189, 191, 190, 190, 180, 169, 147, 138, 136, 136, 139, 139, 143, 139, 140, 145, 151, 157, 156, 159, 151, 155, 140, 141, 131, 138, 134, 140, 141, 146, 147, 146, 147, 150, 153, 146, 147, 154, 146, 153, 153, 155, 162, 178, 172, 172, 176, 179, 193, 194, 200, 197, 199, 193, 195, 193, 193, 199, 199, 194, 197, 195, 188, 177, 177, 170, 178, 174, 175, 173, 172, 181, 180, 179, 172, 176, 173, 174, 177, 170, 169, 173, 168, 176, 172, 185, 212, 221, 220, 225, 220, 226, 226, 225, 225, 225, 223, 223, 220, 223, 220, 222, 221, 221, 220, 221, 221, 221, 220, 222, 222, 221, 223, 219, 219, 217, 219, 219, 217, 217, 216, 216, 217, 219, 216, 215, 215, 216, 213, 217, 215, 212, 216, 211, 212, 208, 211, 209, 213, 213, 210, 209, 204, 196, 194, 188, 180, 180, 179, 178, 176, 174, 178, 178, 174, 176, 178, 173, 174, 167, 175, 168, 165, 165, 166, 170, 167, 167, 164, 159, 165, 163, 161, 161, 164, 161, 159, 160, 160, 158, 159, 161, 159, 158, 163, 163, 163, 160, 164, 161, 161, 160, 159, 161, 154, 158, 150, 157, 157, 157, 157, 159, 152, 155, 153, 152, 156, 159, 158, 157, 153, 160, 162, 157, 157, 160, 159, 161, 161, 160, 161, 166, 163, 166, 169, 168, 172, 168, 167, 168, 167, 166, 167, 174, 171, 166, 165, 164, 164, 164, 162, 162, 167, 168, 170, 165, 168, 164, 169, 157, 187, 182, 176, 179, 78, 181, 182, 186, 186, 190, 185, 167, 145, 141, 141, 139, 138, 144, 147, 145, 148, 148, 163, 166, 166, 163, 159, 155, 146, 139, 134, 138, 140, 144, 145, 150, 149, 146, 148, 155, 155, 153, 155, 151, 153, 153, 154, 151, 162, 172, 167, 175, 175, 176, 192, 196, 198, 198, 194, 198, 193, 197, 199, 198, 195, 198, 196, 195, 187, 175, 178, 172, 174, 177, 172, 169, 169, 172, 182, 176, 168, 169, 172, 174, 174, 170, 171, 172, 172, 177, 177, 190, 211, 220, 220, 222, 220, 225, 225, 224, 225, 224, 225, 221, 220, 224, 222, 220, 218, 219, 219, 219, 223, 221, 219, 220, 219, 220, 220, 218, 214, 216, 215, 217, 219, 219, 218, 218, 218, 218, 216, 214, 216, 214, 213, 214, 215, 214, 212, 214, 214, 213, 213, 212, 213, 213, 209, 208, 202, 195, 191, 186, 185, 178, 174, 176, 177, 178, 179, 184, 180, 177, 183, 177, 178, 170, 175, 176, 172, 163, 169, 166, 166, 172, 162, 163, 161, 161, 168, 169, 168, 165, 159, 159, 163, 163, 161, 160, 161, 161, 163, 164, 162, 160, 159, 159, 162, 160, 161, 166, 161, 158, 158, 154, 160, 163, 165, 159, 153, 159, 155, 152, 163, 161, 159, 157, 160, 164, 163, 166, 162, 161, 165, 164, 160, 161, 161, 167, 164, 164, 166, 166, 172, 173, 173, 168, 168, 168, 168, 171, 165, 168, 166, 169, 165, 164, 162, 164, 166, 168, 166, 167, 168, 169, 171, 162, 184, 184, 183, 182, 81, 182, 190, 188, 187, 188, 182, 163, 140, 145, 144, 141, 146, 153, 157, 154, 154, 159, 161, 174, 170, 167, 163, 149, 151, 143, 138, 144, 138, 142, 144, 150, 153, 151, 153, 156, 162, 158, 151, 150, 153, 155, 156, 157, 161, 177, 170, 173, 181, 178, 194, 199, 193, 196, 191, 195, 189, 197, 200, 201, 199, 199, 195, 198, 184, 174, 177, 171, 174, 171, 171, 171, 170, 171, 178, 180, 171, 174, 172, 178, 179, 178, 176, 179, 180, 179, 181, 193, 211, 216, 217, 221, 218, 221, 224, 223, 226, 225, 225, 222, 219, 220, 214, 219, 219, 218, 218, 217, 220, 220, 220, 220, 219, 223, 221, 217, 216, 215, 215, 216, 217, 216, 214, 220, 217, 219, 215, 214, 216, 217, 213, 215, 216, 216, 211, 213, 212, 212, 214, 206, 215, 212, 206, 206, 201, 197, 187, 183, 180, 181, 178, 182, 181, 181, 181, 183, 180, 184, 179, 177, 178, 172, 175, 179, 176, 166, 163, 167, 167, 165, 172, 166, 168, 169, 170, 171, 163, 165, 162, 164, 166, 163, 157, 161, 163, 165, 163, 163, 162, 163, 162, 167, 167, 164, 166, 158, 165, 157, 159, 162, 158, 163, 160, 162, 157, 163, 159, 160, 158, 158, 157, 163, 161, 161, 160, 162, 158, 165, 161, 163, 158, 160, 162, 164, 163, 164, 165, 166, 171, 172, 171, 164, 170, 167, 168, 172, 168, 170, 164, 167, 165, 160, 167, 158, 163, 164, 168, 170, 173, 172, 166, 159, 189, 183, 176, 180, 74, 177, 186, 186, 188, 187, 183, 164, 145, 148, 141, 144, 149, 154, 156, 158, 162, 160, 172, 172, 170, 169, 154, 146, 150, 148, 142, 143, 143, 149, 149, 147, 151, 146, 157, 157, 160, 155, 156, 155, 157, 158, 159, 159, 167, 176, 172, 173, 181, 179, 189, 196, 191, 198, 193, 194, 195, 193, 198, 197, 198, 201, 198, 195, 190, 174, 178, 179, 174, 174, 166, 169, 175, 168, 181, 176, 174, 182, 182, 174, 181, 181, 174, 179, 179, 178, 180, 192, 215, 216, 220, 221, 222, 220, 222, 224, 225, 224, 223, 222, 221, 220, 218, 219, 218, 217, 218, 218, 220, 222, 219, 221, 220, 222, 217, 214, 214, 216, 215, 218, 217, 219, 217, 220, 218, 217, 214, 215, 216, 216, 217, 214, 213, 214, 214, 213, 215, 216, 213, 214, 214, 211, 210, 206, 202, 192, 187, 184, 185, 182, 181, 183, 181, 184, 185, 183, 185, 183, 183, 182, 177, 174, 182, 179, 182, 170, 170, 168, 172, 174, 176, 171, 173, 175, 169, 175, 165, 168, 165, 167, 169, 164, 163, 168, 165, 164, 170, 165, 169, 170, 175, 173, 171, 168, 171, 162, 169, 163, 167, 169, 161, 161, 161, 162, 162, 158, 162, 158, 161, 162, 162, 161, 163, 156, 165, 158, 157, 164, 159, 162, 155, 156, 160, 160, 165, 160, 163, 165, 166, 172, 172, 167, 171, 168, 172, 168, 171, 167, 164, 170, 169, 170, 160, 168, 169, 172, 169, 176, 171, 170, 170, 161, 185, 182, 177, 185, 80, 184, 188, 190, 188, 186, 184, 160, 150, 148, 144, 150, 153, 157, 163, 161, 164, 161, 175, 171, 167, 172, 156, 153, 159, 149, 146, 144, 149, 151, 152, 151, 150, 153, 154, 162, 159, 161, 162, 161, 165, 157, 162, 163, 163, 176, 171, 173, 179, 179, 188, 193, 194, 190, 191, 193, 191, 190, 197, 198, 198, 198, 195, 194, 188, 179, 178, 179, 176, 172, 173, 174, 176, 173, 180, 179, 179, 180, 181, 183, 182, 184, 172, 180, 179, 179, 179, 188, 212, 216, 219, 217, 222, 219, 223, 222, 224, 221, 222, 218, 222, 221, 220, 220, 217, 216, 216, 218, 222, 221, 216, 217, 220, 219, 220, 218, 214, 218, 217, 219, 217, 218, 214, 214, 216, 218, 215, 215, 217, 215, 215, 211, 216, 214, 216, 213, 212, 215, 216, 209, 211, 209, 206, 203, 201, 190, 186, 187, 181, 183, 184, 180, 180, 182, 185, 183, 183, 181, 180, 181, 177, 177, 180, 173, 179, 182, 170, 172, 171, 174, 180, 177, 171, 172, 175, 167, 169, 172, 166, 169, 170, 168, 170, 170, 170, 175, 172, 173, 175, 176, 176, 174, 177, 175, 173, 175, 172, 175, 171, 168, 166, 167, 165, 165, 161, 157, 158, 160, 163, 159, 162, 162, 165, 163, 164, 162, 157, 155, 161, 156, 150, 159, 161, 163, 165, 164, 166, 172, 173, 174, 174, 170, 170, 168, 172, 172, 180, 177, 177, 181, 176, 178, 176, 180, 180, 184, 181, 181, 178, 179, 179, 175, 178, 180, 180, 184, 89, 181, 189, 184, 188, 187, 182, 161, 150, 144, 145, 150, 154, 160, 167, 165, 167, 168, 171, 170, 171, 162, 157, 154, 157, 154, 150, 150, 147, 152, 148, 154, 155, 156, 162, 166, 166, 167, 168, 174, 173, 168, 163, 165, 167, 177, 176, 174, 183, 181, 185, 191, 193, 192, 186, 192, 189, 188, 193, 199, 196, 195, 196, 193, 189, 178, 176, 173, 174, 168, 175, 170, 176, 174, 177, 177, 186, 182, 188, 180, 185, 181, 179, 181, 183, 185, 178, 192, 210, 213, 220, 221, 222, 220, 221, 220, 223, 221, 220, 221, 220, 220, 220, 216, 215, 216, 220, 221, 220, 218, 212, 216, 215, 215, 219, 215, 216, 214, 218, 218, 215, 213, 216, 214, 212, 218, 214, 215, 213, 215, 215, 216, 215, 213, 213, 216, 214, 209, 211, 210, 210, 210, 206, 202, 190, 189, 191, 188, 188, 186, 182, 183, 181, 185, 184, 181, 186, 185, 180, 180, 180, 173, 176, 174, 176, 181, 177, 167, 171, 177, 170, 176, 172, 173, 171, 171, 168, 173, 170, 176, 174, 171, 171, 172, 179, 177, 177, 174, 179, 176, 182, 180, 176, 177, 173, 175, 174, 171, 170, 171, 166, 170, 163, 165, 158, 157, 163, 164, 162, 160, 162, 164, 167, 163, 162, 164, 162, 162, 165, 162, 157, 163, 164, 166, 174, 178, 177, 179, 180, 181, 180, 181, 184, 182, 183, 186, 189, 185, 187, 187, 185, 185, 190, 187, 190, 190, 187, 187, 187, 188, 185, 179, 182, 178, 174, 182, 71, 180, 185, 187, 184, 183, 177, 160, 151, 150, 150, 153, 160, 166, 164, 165, 169, 168, 172, 170, 167, 168, 153, 155, 153, 155, 152, 149, 152, 152, 154, 153, 168, 166, 166, 175, 177, 177, 177, 178, 179, 171, 166, 165, 169, 175, 173, 175, 182, 183, 191, 188, 192, 186, 186, 186, 189, 190, 194, 198, 192, 195, 193, 197, 190, 175, 178, 174, 176, 169, 173, 172, 174, 179, 180, 183, 183, 182, 187, 180, 179, 185, 175, 180, 181, 186, 183, 194, 209, 212, 218, 221, 220, 218, 220, 222, 221, 220, 221, 217, 218, 217, 219, 218, 213, 216, 218, 221, 216, 215, 216, 212, 213, 213, 213, 210, 213, 214, 217, 218, 215, 214, 217, 215, 214, 215, 214, 208, 214, 219, 214, 215, 215, 214, 212, 213, 216, 211, 208, 211, 211, 206, 205, 194, 187, 183, 189, 188, 188, 187, 184, 185, 181, 187, 184, 184, 186, 181, 184, 184, 182, 176, 177, 176, 177, 175, 174, 171, 176, 172, 172, 171, 172, 173, 175, 172, 171, 173, 175, 176, 176, 179, 177, 178, 175, 176, 176, 173, 173, 173, 177, 175, 176, 176, 172, 174, 170, 169, 168, 171, 168, 171, 170, 170, 167, 162, 165, 167, 168, 160, 160, 164, 167, 167, 165, 161, 164, 163, 164, 164, 168, 169, 172, 184, 184, 188, 192, 193, 189, 193, 193, 192, 194, 189, 186, 194, 199, 190, 195, 199, 201, 202, 202, 205, 206, 204, 205, 203, 206, 207, 206, 207, 197, 192, 189, 202, 115, 192, 188, 185, 178, 175, 180, 166, 158, 156, 160, 154, 159, 166, 167, 166, 161, 166, 170, 168, 171, 165, 154, 158, 162, 158, 150, 149, 151, 151, 153, 157, 162, 161, 165, 166, 174, 169, 167, 172, 173, 169, 161, 163, 169, 170, 169, 174, 176, 172, 180, 181, 179, 181, 180, 171, 178, 179, 183, 186, 186, 185, 188, 184, 177, 166, 166, 154, 161, 163, 158, 162, 165, 163, 169, 170, 169, 168, 172, 169, 171, 172, 163, 163, 169, 173, 175, 181, 194, 192, 192, 200, 198, 195, 202, 200, 201, 202, 200, 198, 200, 201, 196, 197, 194, 195, 198, 197, 207, 202, 198, 201, 193, 189, 191, 183, 190, 189, 190, 192, 192, 192, 192, 188, 187, 185, 187, 186, 196, 206, 199, 194, 193, 188, 192, 190, 192, 194, 193, 199, 203, 210, 213, 211, 206, 190, 208, 191, 190, 185, 192, 199, 195, 179, 180, 177, 174, 164, 188, 177, 172, 159, 152, 152, 148, 153, 144, 148, 156, 160, 172, 160, 157, 160, 164, 163, 170, 161, 161, 193, 187, 196, 189, 204, 206, 187, 176, 193, 170, 154, 139, 138, 139, 140, 135, 158, 149, 149, 147, 160, 142, 153, 166, 140, 147, 150, 137, 154, 166, 148, 133, 131, 133, 134, 152, 136, 137, 151, 139, 134, 136, 137, 132, 141, 145, 146, 150, 151, 147, 149, 149, 159, 156, 163, 188, 163, 151, 144, 141, 140, 155, 134, 130, 146, 131, 152, 147, 140, 137, 142, 155, 159);

--constant memory:MEM_array:=(144, 160, 144, 146, 153, 155, 149, 151, 153, 154, 135, 148, 140, 142, 133, 148, 147, 144, 142, 147, 138, 144, 144, 143, 150, 137, 124, 143, 141, 128, 124, 144, 122, 124, 139, 131, 127, 119, 118, 133, 136, 135, 146, 144, 144, 143, 142, 144, 143, 149, 143, 132, 141, 135, 137, 126, 136, 131, 128, 131, 130, 110, 168, 128, 125, 124, 122, 121, 114, 110, 123, 145, 129, 124, 144, 127, 129, 128, 138, 130, 128, 124, 118, 117, 114, 122, 125, 118, 126, 131, 134, 138, 138, 135, 139, 151, 152, 139, 129, 153, 147, 141, 126, 131, 116, 105, 110, 112, 112, 125, 112, 139, 136, 142, 141, 141, 145, 144, 153, 151, 150, 129, 148, 143, 163, 151, 148, 159, 149, 152, 148, 152, 147, 153, 139, 139, 111, 184, 152, 139, 133, 111, 126, 143, 173, 160, 124, 153, 129, 103, 181, 167, 140, 146, 144, 146, 154, 148, 137, 153, 139, 149, 149, 143, 156, 157, 154, 143, 156, 149, 151, 133, 150, 150, 153, 144, 150, 150, 146, 142, 141, 149, 172, 156, 157, 152, 158, 156, 147, 147, 146, 152, 150, 146, 147, 151, 164, 142, 152, 154, 149, 149, 138, 94, 100, 153, 150, 171, 148, 129, 140, 139, 131, 126, 119, 137, 141, 149, 138, 157, 160, 147, 147, 163, 157, 158, 149, 151, 155, 147, 177, 169, 163, 162, 171, 174, 143, 155, 220, 164, 163, 160, 146, 149, 148, 122, 100, 72, 56, 62, 58, 73, 69, 73, 71, 76, 144, 160, 144, 146, 153, 155, 149, 151, 153, 154, 135, 148, 140, 142, 133, 148, 147, 144, 142, 147, 138, 144, 144, 143, 150, 137, 124, 143, 141, 128, 124, 144, 122, 124, 139, 131, 127, 119, 118, 133, 136, 135, 146, 144, 144, 143, 142, 144, 143, 149, 143, 132, 141, 135, 137, 126, 136, 131, 128, 131, 130, 110, 168, 128, 125, 124, 122, 121, 114, 110, 123, 145, 129, 124, 144, 127, 129, 128, 138, 130, 128, 124, 118, 117, 114, 122, 125, 118, 126, 131, 134, 138, 138, 135, 139, 151, 152, 139, 129, 153, 147, 141, 126, 131, 116, 105, 110, 112, 112, 125, 112, 139, 136, 142, 141, 141, 145, 144, 153, 151, 150, 129, 148, 143, 163, 151, 148, 159, 149, 152, 148, 152, 147, 153, 139, 139, 111, 184, 152, 139, 133, 111, 126, 143, 173, 160, 124, 153, 129, 103, 181, 167, 140, 146, 144, 146, 154, 148, 137, 153, 139, 149, 149, 143, 156, 157, 154, 143, 156, 149, 151, 133, 150, 150, 153, 144, 150, 150, 146, 142, 141, 149, 172, 156, 157, 152, 158, 156, 147, 147, 146, 152, 150, 146, 147, 151, 164, 142, 152, 154, 149, 149, 138, 94, 100, 153, 150, 171, 148, 129, 140, 139, 131, 126, 119, 137, 141, 149, 138, 157, 160, 147, 147, 163, 157, 158, 149, 151, 155, 147, 177, 169, 163, 162, 171, 174, 143, 155, 220, 164, 163, 160, 146, 149, 148, 122, 100, 72, 56, 62, 58, 73, 69, 73, 71, 76, 142, 151, 144, 146, 153, 151, 148, 148, 142, 149, 124, 146, 157, 139, 114, 140, 137, 144, 132, 146, 148, 140, 138, 151, 149, 148, 137, 141, 142, 115, 156, 118, 126, 113, 127, 128, 127, 115, 127, 132, 127, 127, 136, 138, 133, 156, 137, 144, 142, 139, 147, 142, 118, 117, 144, 137, 136, 139, 142, 131, 140, 111, 142, 125, 134, 136, 134, 113, 119, 97, 127, 134, 117, 155, 111, 114, 121, 131, 140, 143, 134, 135, 123, 130, 137, 119, 140, 127, 115, 137, 138, 130, 129, 136, 141, 142, 158, 136, 122, 147, 147, 129, 136, 128, 144, 120, 133, 118, 113, 126, 124, 129, 144, 133, 134, 133, 148, 158, 148, 147, 151, 148, 143, 151, 151, 159, 156, 141, 154, 162, 148, 136, 152, 159, 144, 153, 150, 141, 132, 183, 118, 85, 118, 159, 190, 159, 126, 135, 147, 115, 154, 150, 138, 133, 138, 142, 124, 152, 155, 155, 155, 150, 141, 138, 154, 147, 156, 152, 147, 137, 171, 162, 145, 152, 149, 141, 146, 150, 149, 143, 138, 124, 151, 154, 149, 170, 154, 146, 153, 153, 151, 157, 148, 155, 156, 156, 153, 144, 144, 148, 154, 156, 149, 101, 89, 143, 148, 148, 112, 126, 130, 136, 134, 123, 120, 129, 138, 141, 152, 147, 146, 139, 163, 155, 151, 157, 139, 162, 136, 147, 168, 156, 152, 159, 174, 177, 143, 173, 209, 167, 178, 164, 159, 151, 135, 118, 96, 89, 73, 76, 69, 69, 67, 67, 66, 78, 160, 158, 148, 144, 140, 129, 140, 153, 144, 140, 127, 146, 135, 129, 127, 134, 151, 140, 148, 148, 143, 127, 144, 155, 141, 142, 138, 134, 138, 118, 125, 130, 126, 116, 118, 120, 117, 110, 112, 121, 127, 144, 139, 142, 137, 140, 140, 146, 151, 147, 145, 133, 151, 132, 132, 137, 129, 133, 137, 122, 133, 129, 149, 130, 110, 132, 133, 131, 126, 122, 111, 114, 90, 154, 117, 114, 120, 119, 123, 134, 138, 127, 130, 124, 138, 123, 140, 138, 116, 132, 130, 131, 134, 148, 143, 120, 156, 164, 130, 147, 135, 130, 129, 140, 139, 127, 126, 130, 123, 125, 132, 127, 133, 128, 137, 121, 136, 144, 143, 135, 145, 147, 139, 152, 149, 157, 150, 148, 158, 145, 153, 149, 148, 149, 150, 137, 135, 144, 116, 153, 110, 76, 123, 155, 160, 141, 136, 145, 147, 153, 149, 144, 151, 136, 151, 146, 146, 157, 148, 146, 163, 140, 147, 147, 158, 154, 144, 159, 154, 139, 150, 153, 152, 143, 149, 143, 157, 155, 139, 140, 144, 153, 152, 146, 135, 154, 164, 154, 155, 145, 150, 151, 151, 140, 160, 156, 156, 152, 149, 150, 149, 151, 156, 147, 125, 116, 124, 126, 125, 127, 129, 137, 127, 132, 130, 133, 140, 139, 132, 137, 141, 141, 146, 144, 146, 142, 140, 153, 148, 150, 160, 162, 133, 161, 162, 175, 178, 186, 186, 182, 174, 155, 157, 149, 140, 122, 113, 93, 73, 82, 75, 69, 66, 73, 69, 84, 162, 148, 140, 155, 138, 144, 132, 155, 157, 140, 148, 149, 137, 157, 138, 142, 144, 138, 140, 141, 148, 142, 152, 139, 150, 139, 138, 131, 133, 119, 127, 127, 99, 106, 118, 130, 117, 116, 112, 116, 110, 111, 141, 136, 148, 138, 138, 137, 147, 145, 146, 149, 138, 151, 139, 134, 118, 133, 128, 138, 132, 138, 137, 139, 127, 122, 125, 140, 117, 122, 121, 130, 116, 128, 119, 123, 113, 128, 121, 136, 122, 130, 126, 139, 129, 132, 128, 132, 139, 131, 136, 138, 132, 143, 133, 138, 137, 136, 122, 132, 131, 126, 137, 135, 142, 134, 130, 121, 118, 121, 121, 121, 140, 132, 150, 139, 137, 144, 147, 150, 144, 137, 142, 148, 162, 152, 148, 150, 149, 150, 139, 139, 148, 138, 149, 143, 131, 140, 158, 127, 108, 81, 117, 134, 137, 127, 135, 144, 138, 145, 142, 156, 153, 142, 152, 148, 156, 142, 163, 148, 148, 131, 145, 127, 157, 158, 159, 143, 154, 154, 151, 163, 154, 159, 139, 164, 153, 150, 149, 147, 134, 127, 147, 147, 151, 155, 148, 147, 138, 143, 147, 155, 150, 152, 152, 159, 142, 142, 153, 147, 148, 143, 146, 151, 143, 130, 121, 128, 132, 118, 120, 118, 127, 126, 125, 125, 134, 108, 117, 146, 137, 131, 138, 151, 148, 141, 160, 131, 142, 153, 155, 149, 127, 138, 140, 175, 185, 188, 180, 182, 165, 160, 153, 157, 149, 139, 110, 118, 76, 69, 80, 73, 66, 64, 76, 71, 164, 168, 155, 148, 148, 155, 155, 158, 151, 138, 137, 157, 156, 135, 142, 142, 142, 146, 146, 139, 146, 146, 149, 148, 139, 138, 120, 126, 126, 126, 111, 115, 122, 113, 109, 114, 112, 117, 100, 98, 105, 111, 120, 125, 124, 136, 137, 153, 139, 144, 155, 141, 147, 142, 129, 129, 131, 136, 123, 126, 132, 132, 135, 139, 126, 106, 129, 136, 132, 136, 122, 122, 121, 130, 129, 111, 120, 122, 128, 134, 128, 117, 118, 144, 122, 132, 128, 142, 167, 139, 141, 136, 141, 133, 142, 133, 137, 138, 127, 126, 128, 124, 106, 113, 125, 133, 121, 105, 134, 125, 123, 133, 129, 131, 129, 141, 143, 139, 140, 142, 153, 146, 141, 146, 136, 153, 142, 150, 159, 157, 147, 146, 141, 143, 149, 152, 149, 143, 156, 154, 130, 137, 127, 152, 126, 132, 139, 139, 127, 142, 163, 161, 157, 144, 152, 151, 156, 132, 150, 165, 155, 128, 128, 129, 152, 152, 156, 159, 143, 155, 156, 157, 154, 137, 161, 150, 149, 144, 147, 149, 142, 146, 146, 147, 150, 140, 144, 166, 153, 147, 151, 148, 147, 159, 140, 140, 144, 148, 131, 145, 148, 125, 145, 129, 126, 123, 103, 120, 127, 126, 122, 116, 121, 123, 111, 127, 124, 112, 104, 120, 125, 116, 127, 156, 127, 122, 124, 150, 155, 142, 144, 147, 138, 141, 140, 167, 177, 173, 186, 184, 166, 157, 149, 149, 155, 152, 127, 107, 89, 66, 69, 62, 64, 55, 73, 80, 164, 162, 157, 158, 148, 155, 149, 146, 155, 141, 127, 151, 151, 146, 154, 137, 144, 142, 137, 142, 153, 136, 152, 142, 149, 145, 120, 140, 118, 129, 109, 127, 132, 130, 120, 111, 101, 76, 111, 121, 131, 122, 126, 127, 136, 137, 125, 147, 150, 140, 134, 125, 147, 138, 146, 151, 128, 144, 116, 150, 137, 134, 130, 119, 133, 127, 125, 114, 123, 130, 126, 123, 129, 129, 124, 137, 126, 116, 121, 127, 133, 137, 136, 126, 136, 140, 137, 145, 154, 143, 141, 132, 140, 137, 142, 136, 142, 138, 133, 133, 129, 116, 112, 114, 120, 126, 124, 148, 118, 115, 129, 142, 139, 144, 138, 139, 145, 137, 132, 142, 149, 146, 143, 138, 153, 154, 150, 148, 156, 148, 148, 141, 144, 153, 146, 149, 139, 138, 141, 141, 137, 150, 139, 131, 133, 137, 138, 135, 135, 148, 134, 152, 155, 145, 146, 159, 152, 152, 144, 141, 148, 149, 146, 149, 152, 169, 157, 143, 160, 151, 167, 156, 155, 98, 150, 148, 129, 142, 147, 136, 136, 147, 141, 148, 150, 146, 119, 157, 152, 138, 147, 134, 150, 150, 140, 145, 145, 143, 146, 139, 131, 122, 157, 167, 127, 125, 104, 118, 123, 128, 121, 127, 123, 117, 126, 91, 119, 115, 116, 118, 103, 113, 124, 137, 141, 137, 129, 118, 151, 148, 156, 144, 147, 138, 138, 165, 169, 166, 171, 178, 155, 146, 156, 151, 138, 144, 142, 113, 67, 64, 75, 56, 44, 42, 58, 84, 162, 149, 160, 158, 149, 144, 142, 144, 149, 140, 137, 137, 135, 142, 140, 144, 146, 137, 142, 146, 137, 137, 142, 148, 122, 150, 133, 141, 131, 131, 143, 128, 128, 120, 111, 121, 109, 97, 112, 122, 126, 127, 129, 131, 138, 138, 136, 134, 131, 147, 141, 143, 126, 140, 145, 153, 138, 139, 137, 119, 127, 144, 132, 127, 141, 137, 124, 119, 127, 136, 134, 117, 120, 119, 129, 132, 125, 130, 122, 128, 133, 142, 136, 127, 143, 139, 136, 147, 137, 158, 143, 138, 150, 141, 133, 131, 133, 134, 140, 136, 130, 114, 96, 119, 123, 131, 118, 129, 132, 137, 123, 135, 145, 141, 142, 148, 140, 138, 148, 147, 144, 147, 136, 137, 143, 142, 152, 150, 150, 151, 153, 155, 152, 158, 148, 143, 141, 140, 149, 144, 145, 134, 129, 132, 130, 139, 126, 131, 138, 146, 135, 125, 157, 154, 146, 153, 151, 155, 143, 146, 147, 155, 151, 144, 148, 142, 159, 166, 145, 158, 156, 168, 155, 156, 142, 126, 116, 134, 135, 122, 124, 131, 139, 134, 137, 135, 135, 137, 139, 137, 159, 147, 155, 142, 138, 145, 140, 141, 151, 142, 110, 101, 142, 185, 131, 120, 96, 106, 134, 128, 120, 120, 134, 131, 122, 103, 102, 104, 109, 129, 128, 138, 143, 121, 130, 137, 127, 128, 143, 126, 155, 133, 136, 134, 140, 164, 160, 158, 173, 155, 145, 144, 148, 155, 135, 120, 113, 75, 56, 55, 86, 104, 88, 49, 69, 78, 155, 149, 146, 146, 155, 153, 151, 160, 151, 137, 118, 149, 144, 148, 144, 142, 140, 146, 137, 142, 142, 141, 136, 145, 129, 140, 138, 130, 139, 129, 133, 125, 114, 120, 121, 110, 112, 114, 115, 125, 124, 128, 112, 144, 139, 138, 138, 135, 145, 143, 134, 141, 142, 131, 124, 138, 136, 140, 132, 129, 128, 137, 136, 134, 129, 133, 136, 130, 127, 125, 122, 126, 112, 121, 125, 127, 128, 125, 123, 131, 126, 131, 134, 128, 141, 141, 139, 148, 130, 141, 145, 146, 150, 127, 148, 141, 144, 131, 133, 134, 130, 130, 125, 125, 127, 129, 122, 128, 122, 131, 143, 150, 142, 133, 146, 147, 136, 148, 144, 137, 144, 144, 132, 135, 140, 148, 149, 145, 148, 146, 148, 139, 146, 137, 152, 148, 139, 141, 139, 141, 135, 131, 125, 141, 120, 115, 133, 119, 134, 138, 136, 121, 119, 151, 156, 145, 153, 150, 141, 137, 140, 147, 144, 145, 156, 158, 149, 141, 167, 151, 150, 151, 147, 142, 143, 108, 113, 143, 138, 131, 137, 130, 128, 124, 120, 130, 123, 137, 147, 145, 151, 153, 146, 145, 135, 134, 143, 144, 140, 138, 138, 102, 115, 135, 124, 107, 115, 118, 122, 123, 124, 117, 111, 145, 118, 129, 103, 123, 116, 111, 118, 135, 151, 128, 130, 134, 139, 141, 127, 144, 152, 145, 141, 140, 135, 149, 150, 150, 162, 149, 146, 145, 147, 138, 142, 142, 90, 46, 42, 57, 86, 144, 155, 70, 64, 86, 153, 155, 144, 149, 138, 153, 157, 149, 149, 138, 137, 160, 149, 142, 145, 137, 130, 138, 129, 140, 142, 140, 137, 104, 90, 123, 126, 136, 133, 135, 129, 138, 119, 126, 128, 119, 126, 120, 116, 121, 130, 129, 143, 135, 143, 149, 144, 137, 143, 138, 137, 132, 135, 138, 130, 147, 137, 130, 132, 139, 133, 142, 129, 133, 130, 138, 126, 136, 128, 120, 122, 129, 127, 127, 123, 134, 127, 123, 128, 132, 130, 123, 140, 130, 142, 144, 127, 129, 144, 141, 138, 142, 141, 138, 135, 128, 135, 129, 133, 143, 138, 130, 133, 136, 140, 123, 122, 112, 133, 134, 133, 142, 132, 165, 137, 148, 138, 149, 144, 153, 143, 139, 149, 144, 155, 143, 143, 155, 149, 143, 145, 150, 141, 141, 136, 133, 137, 136, 135, 144, 143, 138, 137, 120, 168, 119, 127, 130, 132, 119, 145, 134, 143, 137, 134, 138, 153, 142, 147, 142, 134, 152, 144, 143, 144, 147, 149, 150, 148, 152, 153, 149, 155, 141, 147, 143, 130, 146, 122, 142, 137, 133, 119, 128, 128, 126, 116, 126, 120, 151, 149, 149, 150, 127, 179, 128, 132, 141, 133, 133, 128, 126, 131, 116, 107, 93, 109, 121, 121, 116, 131, 124, 121, 138, 125, 138, 127, 124, 123, 109, 114, 122, 140, 128, 138, 126, 155, 128, 124, 152, 180, 159, 156, 145, 144, 146, 140, 148, 151, 143, 137, 142, 144, 148, 155, 155, 86, 5, 18, 46, 84, 177, 175, 114, 75, 111, 160, 158, 153, 146, 151, 158, 144, 149, 144, 140, 155, 144, 140, 138, 148, 148, 136, 137, 112, 110, 144, 138, 146, 120, 119, 131, 123, 129, 131, 133, 118, 132, 127, 127, 125, 109, 116, 132, 130, 132, 133, 133, 137, 140, 137, 142, 146, 137, 136, 139, 128, 130, 136, 126, 132, 151, 137, 132, 136, 135, 134, 133, 128, 140, 131, 131, 128, 129, 115, 118, 130, 130, 133, 116, 121, 129, 131, 123, 150, 128, 126, 128, 127, 137, 136, 136, 132, 137, 127, 143, 137, 136, 140, 138, 135, 141, 145, 122, 128, 168, 138, 136, 128, 137, 148, 139, 131, 132, 131, 131, 133, 123, 103, 137, 134, 141, 149, 149, 145, 137, 129, 150, 142, 131, 152, 154, 140, 153, 145, 148, 141, 134, 137, 136, 130, 139, 140, 138, 128, 135, 129, 118, 142, 121, 155, 131, 133, 108, 128, 110, 125, 139, 132, 133, 142, 152, 144, 145, 137, 176, 146, 141, 147, 157, 142, 146, 135, 134, 137, 170, 153, 149, 141, 138, 144, 136, 147, 141, 129, 146, 145, 112, 131, 155, 128, 125, 92, 153, 156, 148, 149, 143, 142, 137, 147, 131, 133, 137, 136, 127, 119, 127, 118, 104, 87, 121, 110, 122, 110, 130, 130, 134, 123, 124, 135, 134, 135, 131, 119, 108, 117, 118, 111, 137, 133, 150, 141, 115, 118, 140, 172, 189, 156, 181, 151, 137, 136, 148, 144, 144, 135, 140, 144, 131, 148, 172, 99, 15, 12, 25, 90, 177, 184, 137, 100, 126, 160, 158, 157, 133, 149, 171, 146, 149, 140, 140, 152, 144, 144, 146, 135, 146, 142, 137, 133, 122, 132, 142, 138, 139, 127, 128, 119, 129, 138, 141, 133, 131, 125, 119, 136, 132, 131, 124, 140, 142, 141, 135, 138, 139, 141, 146, 140, 145, 140, 135, 141, 126, 131, 134, 144, 139, 141, 125, 123, 123, 121, 137, 124, 142, 128, 132, 115, 151, 108, 124, 134, 124, 123, 119, 115, 126, 126, 120, 133, 131, 125, 131, 126, 126, 120, 137, 131, 131, 135, 145, 141, 142, 134, 134, 134, 134, 139, 132, 135, 129, 130, 136, 143, 125, 141, 137, 134, 137, 134, 126, 127, 131, 136, 142, 137, 136, 138, 128, 132, 144, 139, 136, 141, 139, 148, 139, 138, 138, 149, 149, 150, 152, 142, 145, 144, 139, 144, 137, 139, 142, 126, 136, 119, 129, 133, 122, 126, 133, 126, 132, 127, 136, 141, 148, 143, 150, 159, 156, 138, 159, 141, 146, 143, 159, 146, 144, 150, 147, 154, 152, 153, 135, 142, 139, 139, 147, 141, 141, 130, 134, 130, 93, 118, 174, 128, 124, 88, 134, 170, 142, 147, 148, 147, 145, 138, 139, 132, 129, 140, 130, 131, 133, 129, 127, 113, 100, 107, 125, 120, 127, 136, 137, 123, 132, 132, 137, 132, 129, 112, 120, 126, 118, 114, 151, 137, 154, 149, 109, 110, 134, 161, 174, 141, 174, 165, 157, 142, 138, 125, 154, 160, 134, 141, 138, 150, 153, 120, 18, 0, 28, 94, 154, 177, 125, 115, 152, 155, 155, 148, 132, 157, 161, 143, 149, 151, 139, 156, 148, 144, 150, 139, 144, 140, 144, 137, 142, 137, 149, 143, 130, 130, 117, 131, 119, 124, 128, 133, 127, 141, 136, 132, 135, 132, 139, 135, 132, 138, 139, 141, 139, 145, 141, 140, 138, 147, 120, 112, 133, 136, 139, 154, 133, 129, 132, 149, 138, 129, 132, 138, 130, 117, 125, 105, 126, 138, 125, 120, 127, 139, 131, 134, 132, 133, 132, 117, 121, 132, 131, 130, 125, 134, 130, 135, 134, 125, 140, 142, 126, 128, 131, 127, 133, 132, 128, 130, 138, 143, 137, 137, 137, 138, 137, 130, 137, 125, 140, 117, 135, 143, 137, 138, 131, 139, 123, 118, 135, 138, 134, 149, 146, 144, 135, 134, 147, 139, 143, 147, 143, 144, 150, 136, 135, 135, 131, 138, 129, 126, 127, 136, 125, 131, 132, 130, 131, 123, 131, 134, 150, 128, 137, 140, 146, 139, 144, 133, 154, 149, 164, 148, 145, 127, 163, 149, 148, 143, 145, 143, 139, 145, 136, 142, 141, 138, 146, 138, 141, 137, 121, 108, 137, 121, 136, 124, 134, 136, 134, 144, 147, 139, 156, 137, 138, 142, 131, 114, 136, 126, 131, 124, 134, 123, 114, 114, 123, 138, 131, 119, 150, 137, 131, 136, 140, 119, 117, 123, 123, 128, 124, 108, 157, 139, 140, 174, 145, 130, 132, 151, 157, 156, 156, 155, 155, 155, 107, 69, 180, 226, 123, 129, 142, 127, 154, 158, 81, 18, 20, 70, 123, 136, 129, 123, 182, 143, 153, 149, 144, 151, 151, 149, 146, 144, 151, 151, 148, 146, 143, 152, 144, 146, 143, 132, 140, 136, 148, 134, 120, 129, 141, 136, 108, 115, 143, 140, 125, 138, 138, 133, 124, 132, 154, 148, 139, 138, 141, 135, 143, 130, 146, 145, 149, 144, 140, 126, 130, 124, 134, 135, 137, 137, 134, 136, 134, 131, 132, 128, 131, 120, 125, 126, 127, 127, 123, 115, 126, 120, 124, 141, 131, 135, 133, 133, 136, 132, 135, 130, 130, 134, 127, 135, 137, 126, 139, 132, 121, 126, 123, 130, 123, 134, 123, 137, 142, 133, 129, 142, 139, 140, 134, 126, 131, 121, 131, 129, 127, 136, 143, 135, 135, 138, 139, 128, 139, 130, 132, 139, 136, 137, 150, 149, 136, 138, 144, 134, 132, 135, 140, 131, 136, 145, 128, 142, 127, 112, 105, 138, 134, 120, 122, 134, 127, 133, 135, 141, 137, 144, 148, 171, 151, 157, 145, 166, 145, 134, 151, 141, 137, 139, 148, 132, 147, 168, 142, 146, 144, 127, 133, 136, 141, 144, 146, 141, 152, 161, 130, 127, 121, 112, 133, 142, 151, 130, 149, 152, 154, 151, 151, 143, 142, 133, 142, 127, 122, 130, 124, 134, 136, 112, 111, 116, 114, 115, 124, 132, 117, 132, 138, 138, 147, 126, 98, 167, 138, 130, 127, 132, 146, 142, 146, 154, 141, 172, 146, 142, 149, 148, 164, 162, 152, 159, 92, 39, 145, 206, 123, 132, 129, 131, 133, 154, 124, 78, 34, 51, 92, 100, 120, 153, 182, 149, 151, 157, 149, 152, 146, 155, 144, 141, 146, 153, 151, 152, 144, 140, 141, 140, 142, 136, 148, 133, 122, 97, 98, 134, 191, 211, 145, 113, 117, 145, 141, 142, 144, 138, 144, 137, 140, 139, 151, 131, 133, 138, 145, 143, 134, 147, 135, 137, 133, 136, 135, 130, 137, 130, 132, 140, 126, 138, 135, 139, 112, 115, 119, 119, 132, 138, 132, 138, 136, 132, 127, 138, 136, 127, 135, 139, 119, 132, 139, 122, 127, 130, 136, 128, 127, 131, 131, 139, 129, 129, 137, 132, 126, 136, 133, 123, 126, 139, 141, 129, 133, 127, 146, 134, 131, 130, 130, 128, 126, 126, 124, 143, 129, 117, 143, 132, 139, 141, 119, 138, 138, 133, 128, 142, 140, 148, 146, 138, 142, 130, 140, 133, 139, 138, 135, 147, 135, 132, 127, 121, 117, 123, 115, 136, 126, 126, 127, 119, 137, 139, 134, 145, 149, 136, 128, 163, 173, 152, 151, 147, 148, 140, 143, 145, 150, 115, 139, 162, 140, 142, 147, 141, 133, 140, 141, 144, 147, 142, 145, 144, 144, 133, 128, 119, 121, 130, 168, 144, 150, 149, 153, 156, 138, 139, 133, 135, 143, 139, 134, 132, 132, 127, 131, 145, 125, 129, 118, 131, 121, 135, 130, 128, 141, 140, 142, 144, 115, 146, 141, 145, 143, 135, 145, 147, 156, 159, 132, 155, 165, 139, 143, 139, 148, 157, 157, 156, 136, 79, 115, 136, 119, 127, 131, 132, 139, 146, 148, 104, 77, 67, 80, 93, 120, 164, 196, 149, 148, 157, 146, 148, 155, 153, 151, 149, 149, 149, 144, 144, 141, 129, 140, 144, 145, 152, 149, 130, 92, 66, 82, 127, 189, 234, 225, 134, 108, 135, 130, 146, 138, 141, 143, 140, 141, 141, 139, 137, 137, 147, 139, 140, 139, 135, 148, 147, 137, 142, 141, 130, 126, 116, 128, 131, 124, 135, 137, 136, 127, 121, 124, 133, 130, 129, 133, 123, 118, 147, 129, 145, 132, 132, 133, 136, 129, 120, 118, 128, 131, 129, 130, 135, 134, 133, 127, 128, 121, 132, 131, 133, 143, 138, 151, 129, 125, 149, 145, 135, 133, 136, 128, 129, 118, 125, 128, 119, 128, 131, 142, 139, 134, 132, 129, 133, 134, 134, 126, 126, 142, 127, 131, 132, 149, 134, 137, 137, 134, 129, 142, 131, 134, 145, 141, 132, 141, 127, 137, 120, 132, 122, 118, 130, 132, 124, 130, 120, 137, 141, 140, 142, 147, 130, 125, 156, 173, 145, 147, 143, 151, 139, 134, 152, 152, 139, 139, 139, 136, 136, 141, 137, 143, 132, 138, 138, 151, 136, 137, 142, 140, 135, 140, 128, 126, 134, 152, 131, 138, 141, 146, 142, 138, 145, 137, 129, 132, 132, 127, 117, 138, 142, 130, 135, 123, 127, 127, 132, 128, 129, 140, 142, 147, 146, 154, 182, 151, 144, 148, 148, 144, 151, 143, 144, 153, 156, 135, 141, 141, 138, 149, 149, 152, 161, 148, 141, 131, 130, 132, 131, 137, 132, 130, 127, 135, 147, 135, 96, 94, 89, 97, 104, 131, 163, 173, 153, 155, 146, 131, 138, 155, 161, 151, 153, 147, 136, 149, 139, 132, 140, 149, 148, 156, 159, 158, 125, 56, 42, 59, 112, 181, 238, 240, 186, 110, 133, 133, 142, 147, 139, 134, 141, 148, 144, 143, 147, 145, 144, 148, 140, 145, 128, 120, 137, 137, 139, 135, 141, 131, 134, 127, 129, 125, 134, 131, 137, 121, 92, 121, 139, 150, 132, 135, 115, 119, 132, 132, 127, 129, 136, 121, 135, 126, 117, 130, 130, 121, 137, 130, 132, 127, 130, 133, 129, 119, 140, 137, 127, 138, 131, 134, 139, 126, 142, 153, 146, 133, 135, 133, 138, 143, 134, 131, 132, 126, 131, 140, 142, 143, 133, 135, 139, 143, 146, 121, 146, 133, 123, 119, 159, 184, 142, 136, 136, 135, 139, 129, 142, 142, 137, 144, 134, 140, 142, 133, 132, 132, 129, 130, 120, 146, 135, 133, 141, 153, 147, 120, 157, 148, 151, 124, 147, 153, 140, 152, 157, 151, 152, 150, 140, 140, 128, 155, 151, 150, 138, 143, 137, 148, 143, 130, 137, 150, 143, 134, 137, 148, 141, 135, 143, 140, 133, 131, 110, 149, 149, 134, 143, 135, 138, 128, 131, 128, 126, 133, 124, 128, 136, 140, 126, 133, 132, 124, 145, 113, 139, 141, 141, 149, 153, 150, 133, 166, 152, 156, 148, 138, 145, 150, 156, 154, 156, 158, 147, 143, 146, 157, 155, 157, 150, 141, 136, 133, 142, 130, 137, 144, 138, 137, 135, 133, 127, 131, 110, 86, 95, 107, 109, 121, 135, 174, 157, 158, 142, 136, 149, 147, 155, 149, 148, 152, 139, 155, 148, 146, 146, 144, 147, 140, 157, 171, 123, 51, 29, 54, 107, 127, 228, 236, 192, 103, 115, 147, 137, 145, 133, 146, 148, 125, 159, 144, 139, 143, 149, 146, 147, 141, 140, 137, 139, 143, 129, 136, 127, 129, 133, 133, 141, 135, 132, 134, 114, 136, 151, 136, 120, 127, 142, 133, 137, 131, 140, 130, 143, 128, 128, 125, 135, 126, 117, 130, 130, 131, 134, 136, 137, 129, 124, 123, 134, 129, 126, 138, 134, 145, 137, 140, 143, 136, 123, 143, 142, 135, 143, 139, 142, 150, 146, 136, 137, 128, 125, 108, 150, 163, 133, 124, 141, 137, 138, 132, 123, 133, 107, 102, 150, 176, 148, 126, 140, 133, 133, 135, 138, 146, 136, 137, 132, 136, 133, 135, 134, 140, 132, 138, 124, 138, 148, 145, 134, 145, 148, 154, 146, 146, 149, 141, 145, 146, 147, 142, 139, 150, 153, 152, 131, 166, 143, 145, 144, 144, 153, 140, 139, 138, 143, 141, 146, 140, 149, 155, 149, 139, 154, 141, 138, 152, 146, 146, 134, 131, 136, 134, 142, 137, 131, 134, 130, 132, 142, 131, 133, 145, 128, 135, 124, 140, 131, 126, 141, 132, 130, 141, 138, 138, 142, 155, 135, 153, 151, 139, 146, 147, 128, 148, 145, 150, 154, 155, 152, 157, 153, 148, 152, 156, 154, 145, 132, 138, 137, 131, 142, 142, 140, 127, 126, 131, 138, 133, 123, 98, 102, 111, 120, 117, 153, 157, 149, 148, 145, 143, 148, 155, 151, 153, 155, 149, 153, 144, 144, 143, 148, 141, 147, 144, 149, 157, 139, 45, 19, 48, 85, 121, 190, 222, 157, 110, 121, 131, 137, 136, 140, 139, 143, 145, 141, 133, 132, 143, 139, 141, 138, 137, 139, 134, 134, 121, 138, 143, 139, 137, 129, 135, 130, 130, 138, 132, 112, 119, 125, 167, 129, 141, 125, 133, 135, 127, 132, 114, 126, 125, 127, 126, 123, 114, 114, 123, 120, 123, 129, 124, 135, 133, 130, 124, 126, 132, 137, 131, 132, 134, 127, 143, 139, 136, 143, 125, 136, 125, 146, 147, 135, 141, 137, 134, 135, 137, 135, 115, 137, 152, 123, 135, 135, 144, 131, 133, 136, 137, 130, 105, 139, 145, 136, 129, 140, 135, 140, 141, 139, 137, 146, 131, 137, 134, 133, 126, 129, 126, 139, 132, 154, 151, 145, 153, 143, 145, 141, 153, 158, 153, 141, 143, 145, 149, 155, 154, 148, 152, 149, 155, 150, 141, 142, 146, 147, 144, 155, 138, 146, 140, 133, 128, 143, 142, 149, 149, 147, 153, 142, 149, 140, 134, 137, 132, 138, 142, 135, 130, 134, 131, 139, 137, 140, 128, 129, 125, 127, 146, 125, 130, 137, 128, 141, 135, 125, 135, 132, 144, 146, 143, 160, 143, 148, 144, 141, 143, 149, 146, 154, 130, 149, 154, 151, 148, 154, 156, 141, 143, 148, 153, 155, 151, 143, 146, 135, 143, 148, 140, 140, 128, 124, 119, 129, 142, 127, 119, 99, 106, 118, 135, 138, 161, 155, 143, 153, 151, 150, 159, 151, 143, 146, 146, 144, 148, 150, 142, 144, 146, 134, 138, 149, 155, 148, 91, 34, 40, 68, 111, 154, 138, 140, 118, 133, 137, 131, 136, 148, 148, 137, 137, 143, 140, 136, 127, 138, 136, 127, 144, 128, 133, 126, 127, 130, 137, 139, 133, 125, 123, 144, 134, 138, 148, 145, 141, 117, 153, 128, 134, 133, 124, 134, 129, 125, 133, 130, 127, 130, 125, 126, 100, 89, 118, 123, 120, 117, 121, 116, 143, 127, 133, 130, 129, 131, 128, 148, 140, 136, 139, 139, 141, 138, 145, 124, 121, 138, 144, 137, 140, 141, 135, 133, 127, 139, 141, 142, 146, 129, 132, 148, 145, 128, 128, 151, 130, 130, 115, 128, 128, 126, 126, 137, 145, 131, 136, 138, 142, 130, 141, 140, 119, 135, 131, 132, 133, 137, 131, 148, 146, 148, 152, 152, 145, 150, 151, 146, 144, 139, 140, 140, 146, 150, 145, 160, 147, 153, 143, 149, 139, 146, 146, 150, 143, 149, 135, 133, 126, 143, 135, 140, 150, 138, 162, 162, 154, 155, 141, 144, 142, 128, 143, 130, 128, 111, 124, 115, 112, 135, 137, 137, 129, 132, 130, 139, 135, 130, 133, 133, 130, 138, 131, 126, 117, 129, 136, 138, 152, 144, 128, 149, 141, 140, 140, 142, 137, 145, 138, 146, 149, 147, 144, 146, 151, 143, 154, 151, 154, 144, 148, 146, 148, 133, 143, 146, 138, 137, 137, 121, 141, 124, 138, 144, 130, 129, 115, 108, 127, 142, 169, 158, 164, 147, 145, 154, 151, 152, 140, 148, 151, 149, 145, 132, 148, 151, 150, 139, 142, 145, 155, 148, 145, 110, 68, 89, 110, 116, 127, 135, 144, 141, 134, 142, 141, 139, 134, 147, 134, 140, 137, 147, 137, 141, 130, 138, 133, 135, 139, 136, 138, 130, 127, 133, 117, 119, 139, 155, 142, 132, 139, 131, 140, 136, 141, 128, 138, 136, 141, 143, 132, 132, 133, 120, 129, 124, 118, 114, 97, 120, 130, 134, 117, 123, 130, 136, 136, 130, 129, 134, 122, 128, 127, 134, 130, 132, 140, 136, 135, 149, 132, 134, 127, 129, 141, 135, 150, 149, 133, 142, 137, 140, 128, 144, 137, 145, 135, 140, 143, 109, 121, 129, 119, 137, 140, 138, 136, 134, 130, 129, 137, 132, 143, 135, 136, 140, 133, 142, 139, 133, 131, 139, 147, 142, 138, 148, 138, 156, 149, 151, 141, 147, 144, 157, 155, 148, 147, 149, 153, 147, 153, 156, 144, 145, 152, 159, 153, 145, 147, 145, 136, 151, 144, 149, 143, 147, 146, 145, 146, 150, 151, 131, 150, 173, 148, 137, 126, 134, 147, 136, 136, 139, 124, 125, 128, 136, 139, 133, 134, 145, 134, 125, 150, 144, 139, 132, 151, 131, 128, 128, 128, 131, 136, 131, 137, 146, 135, 138, 142, 137, 137, 127, 132, 137, 137, 137, 149, 149, 152, 148, 153, 152, 151, 149, 145, 146, 146, 144, 148, 139, 141, 149, 140, 135, 137, 146, 135, 129, 135, 140, 127, 126, 119, 101, 115, 144, 158, 158, 150, 139, 149, 158, 155, 148, 148, 149, 146, 152, 149, 135, 140, 150, 141, 149, 148, 147, 152, 139, 145, 152, 142, 140, 118, 122, 136, 148, 154, 146, 138, 139, 138, 145, 134, 144, 148, 146, 137, 149, 141, 133, 137, 133, 132, 145, 144, 116, 160, 126, 128, 126, 118, 114, 127, 158, 137, 132, 136, 119, 136, 139, 124, 175, 132, 133, 136, 133, 132, 136, 132, 120, 126, 130, 133, 126, 127, 122, 124, 120, 141, 126, 129, 133, 139, 132, 136, 129, 123, 153, 126, 131, 141, 138, 137, 139, 147, 136, 134, 139, 146, 139, 139, 131, 137, 129, 132, 129, 145, 141, 136, 144, 141, 146, 131, 132, 138, 108, 135, 155, 140, 124, 133, 122, 136, 124, 126, 124, 137, 132, 141, 137, 136, 131, 129, 128, 142, 142, 142, 142, 143, 145, 149, 152, 149, 147, 149, 143, 150, 154, 151, 157, 145, 148, 140, 148, 157, 139, 132, 175, 156, 148, 146, 151, 153, 143, 145, 141, 130, 147, 142, 141, 138, 148, 149, 156, 142, 157, 149, 142, 136, 146, 154, 146, 140, 150, 155, 141, 137, 138, 133, 130, 140, 138, 145, 131, 135, 142, 141, 140, 133, 138, 139, 127, 136, 138, 134, 136, 140, 129, 126, 146, 145, 140, 137, 135, 137, 132, 128, 116, 119, 128, 131, 123, 149, 151, 145, 143, 139, 152, 158, 154, 143, 148, 146, 146, 154, 140, 143, 148, 140, 132, 142, 144, 137, 144, 135, 142, 137, 143, 141, 112, 118, 131, 158, 152, 163, 154, 148, 148, 148, 143, 144, 142, 148, 151, 147, 142, 142, 153, 149, 144, 149, 150, 157, 157, 149, 153, 144, 145, 141, 134, 137, 144, 138, 146, 129, 141, 144, 141, 150, 139, 144, 146, 138, 148, 145, 132, 133, 129, 138, 142, 144, 144, 131, 127, 134, 113, 119, 119, 152, 155, 144, 138, 131, 132, 136, 124, 108, 145, 131, 137, 141, 134, 147, 135, 108, 117, 127, 127, 138, 131, 129, 126, 118, 125, 122, 129, 127, 135, 132, 134, 134, 125, 124, 132, 124, 131, 143, 144, 138, 137, 146, 135, 140, 140, 136, 140, 147, 137, 145, 149, 120, 130, 134, 133, 143, 142, 126, 110, 169, 140, 133, 98, 125, 159, 174, 133, 132, 129, 132, 125, 129, 133, 134, 133, 141, 138, 125, 133, 132, 141, 133, 140, 150, 137, 143, 151, 143, 146, 151, 151, 149, 146, 150, 152, 146, 152, 142, 145, 155, 148, 154, 147, 149, 139, 150, 146, 151, 156, 140, 147, 153, 134, 141, 145, 143, 144, 147, 152, 140, 154, 146, 149, 148, 152, 148, 142, 144, 144, 141, 144, 145, 139, 137, 143, 138, 124, 131, 136, 137, 135, 136, 122, 141, 163, 138, 130, 141, 130, 124, 139, 142, 140, 135, 153, 144, 134, 140, 144, 147, 138, 141, 135, 128, 123, 126, 115, 129, 117, 132, 157, 149, 141, 141, 146, 152, 155, 143, 150, 148, 143, 139, 156, 130, 144, 137, 148, 146, 147, 144, 129, 128, 143, 137, 140, 153, 129, 116, 126, 140, 156, 153, 143, 139, 146, 135, 138, 138, 149, 144, 148, 143, 156, 146, 148, 149, 150, 144, 152, 150, 144, 144, 152, 144, 143, 145, 144, 142, 138, 140, 137, 137, 144, 141, 144, 145, 142, 139, 140, 140, 138, 134, 136, 135, 138, 137, 130, 148, 142, 137, 127, 145, 159, 131, 125, 133, 146, 143, 139, 136, 136, 130, 131, 131, 125, 133, 134, 124, 130, 138, 137, 135, 124, 131, 127, 133, 131, 135, 124, 112, 133, 129, 126, 129, 137, 135, 132, 131, 134, 127, 137, 120, 128, 140, 135, 134, 136, 135, 142, 144, 139, 129, 134, 133, 118, 156, 167, 145, 134, 129, 130, 146, 135, 141, 125, 144, 145, 126, 91, 117, 153, 155, 120, 131, 132, 145, 127, 127, 128, 127, 132, 136, 134, 139, 142, 139, 132, 141, 142, 142, 137, 148, 141, 141, 151, 155, 154, 144, 141, 149, 152, 149, 154, 152, 153, 154, 145, 145, 146, 145, 147, 148, 149, 153, 146, 144, 144, 157, 132, 153, 158, 152, 132, 151, 141, 151, 161, 155, 138, 148, 146, 153, 145, 134, 141, 150, 145, 152, 140, 144, 149, 149, 144, 138, 146, 134, 146, 148, 135, 135, 152, 141, 132, 124, 130, 137, 136, 148, 152, 152, 150, 147, 137, 143, 159, 156, 130, 133, 124, 127, 136, 127, 124, 118, 112, 145, 147, 143, 149, 153, 153, 154, 149, 151, 152, 143, 135, 126, 159, 146, 134, 141, 140, 137, 152, 143, 120, 121, 154, 137, 146, 153, 134, 141, 128, 138, 144, 156, 132, 130, 166, 153, 144, 144, 151, 148, 151, 148, 149, 141, 153, 150, 151, 145, 152, 143, 148, 141, 153, 144, 145, 144, 148, 142, 137, 134, 144, 142, 139, 141, 133, 138, 143, 133, 141, 127, 130, 138, 137, 138, 138, 140, 134, 132, 136, 133, 104, 134, 151, 141, 124, 129, 145, 137, 135, 135, 130, 132, 137, 136, 121, 172, 156, 126, 123, 131, 131, 133, 130, 127, 132, 136, 129, 133, 123, 118, 121, 124, 133, 133, 131, 114, 162, 143, 120, 129, 135, 138, 123, 138, 135, 137, 137, 132, 133, 132, 149, 138, 140, 133, 120, 145, 160, 138, 139, 132, 134, 146, 139, 133, 138, 137, 138, 137, 128, 113, 134, 129, 117, 128, 130, 134, 134, 123, 129, 124, 122, 135, 133, 126, 140, 134, 141, 147, 137, 149, 137, 142, 156, 150, 145, 146, 148, 154, 146, 148, 157, 145, 148, 152, 142, 152, 160, 165, 141, 145, 147, 153, 149, 149, 150, 147, 145, 138, 135, 160, 158, 153, 151, 152, 145, 147, 156, 151, 160, 151, 144, 136, 150, 147, 141, 148, 148, 146, 151, 142, 154, 146, 140, 147, 130, 133, 133, 151, 149, 151, 138, 145, 140, 140, 134, 141, 143, 145, 150, 154, 146, 150, 143, 128, 153, 155, 129, 137, 123, 127, 131, 119, 123, 122, 121, 127, 135, 147, 148, 152, 158, 161, 149, 148, 149, 151, 154, 145, 153, 148, 143, 137, 151, 149, 148, 154, 137, 121, 149, 140, 145, 140, 151, 157, 149, 141, 147, 149, 105, 121, 168, 199, 139, 134, 148, 149, 148, 157, 144, 154, 147, 143, 149, 151, 149, 152, 156, 156, 143, 150, 142, 136, 142, 144, 140, 140, 144, 144, 142, 125, 131, 140, 135, 138, 133, 137, 131, 140, 142, 144, 140, 137, 137, 127, 136, 130, 132, 137, 129, 127, 128, 123, 121, 117, 121, 126, 115, 129, 135, 109, 96, 137, 169, 122, 129, 137, 132, 128, 125, 122, 130, 130, 136, 138, 125, 115, 120, 128, 124, 127, 121, 88, 135, 149, 135, 132, 129, 134, 132, 135, 133, 139, 134, 141, 137, 139, 138, 130, 133, 144, 130, 135, 139, 132, 145, 132, 142, 150, 140, 138, 146, 134, 129, 121, 157, 123, 131, 118, 116, 125, 122, 133, 136, 138, 137, 135, 132, 120, 128, 133, 105, 129, 127, 137, 149, 149, 145, 152, 152, 150, 151, 147, 154, 146, 149, 149, 140, 147, 155, 146, 133, 150, 174, 197, 165, 148, 148, 157, 151, 148, 148, 149, 152, 146, 143, 150, 148, 143, 148, 148, 138, 135, 150, 146, 157, 151, 159, 151, 137, 154, 143, 138, 135, 145, 155, 147, 151, 150, 142, 139, 149, 137, 130, 147, 153, 144, 142, 139, 146, 146, 141, 141, 148, 146, 159, 158, 155, 144, 148, 132, 147, 141, 139, 138, 139, 133, 127, 126, 131, 116, 119, 131, 135, 138, 144, 149, 157, 151, 154, 150, 154, 148, 147, 158, 145, 140, 148, 146, 157, 147, 158, 146, 133, 142, 146, 140, 136, 138, 156, 155, 146, 148, 131, 139, 94, 99, 154, 176, 147, 140, 139, 145, 153, 151, 153, 145, 148, 147, 141, 153, 152, 152, 148, 141, 132, 146, 144, 143, 147, 142, 146, 144, 142, 142, 145, 135, 134, 140, 121, 140, 146, 135, 141, 151, 140, 132, 147, 144, 123, 129, 138, 141, 131, 141, 121, 121, 135, 139, 130, 125, 133, 123, 127, 127, 136, 126, 100, 119, 125, 121, 125, 128, 130, 127, 118, 130, 122, 125, 133, 132, 134, 129, 126, 128, 105, 110, 125, 117, 110, 120, 132, 136, 135, 137, 131, 132, 143, 142, 137, 138, 145, 133, 146, 137, 141, 140, 139, 140, 140, 116, 138, 146, 137, 139, 137, 141, 136, 138, 138, 123, 128, 123, 135, 137, 128, 127, 126, 109, 136, 127, 126, 135, 129, 127, 140, 140, 129, 135, 128, 142, 142, 147, 151, 155, 144, 137, 138, 149, 135, 150, 152, 142, 161, 144, 143, 122, 118, 143, 163, 188, 167, 157, 152, 151, 155, 142, 156, 146, 149, 156, 156, 152, 151, 149, 153, 150, 151, 150, 147, 150, 150, 150, 151, 139, 149, 143, 148, 143, 144, 125, 153, 154, 144, 151, 149, 137, 148, 138, 143, 140, 141, 150, 136, 137, 145, 150, 147, 137, 162, 153, 147, 160, 162, 148, 154, 151, 140, 145, 137, 148, 145, 127, 133, 127, 127, 120, 120, 127, 133, 138, 151, 152, 153, 156, 147, 148, 157, 154, 152, 151, 143, 147, 149, 151, 150, 159, 168, 147, 140, 138, 149, 142, 146, 150, 147, 152, 156, 142, 156, 142, 128, 113, 136, 150, 140, 146, 141, 150, 146, 154, 145, 154, 148, 141, 149, 159, 149, 147, 154, 147, 143, 143, 147, 142, 144, 147, 146, 148, 142, 142, 137, 130, 133, 133, 135, 146, 140, 139, 143, 147, 137, 133, 140, 139, 136, 125, 130, 139, 138, 144, 141, 131, 130, 134, 138, 117, 124, 131, 132, 125, 119, 101, 93, 117, 124, 117, 109, 134, 130, 123, 124, 133, 128, 119, 119, 136, 133, 117, 121, 124, 116, 116, 124, 130, 124, 113, 119, 123, 123, 126, 135, 139, 141, 134, 134, 135, 135, 144, 134, 145, 137, 139, 133, 133, 138, 137, 132, 131, 141, 135, 128, 137, 134, 135, 139, 129, 131, 133, 129, 133, 142, 137, 122, 101, 140, 144, 129, 140, 133, 119, 142, 141, 131, 138, 130, 141, 137, 151, 152, 147, 144, 151, 150, 152, 150, 147, 137, 143, 146, 146, 148, 140, 106, 136, 147, 179, 161, 138, 145, 135, 165, 151, 152, 143, 152, 153, 157, 152, 151, 157, 143, 148, 154, 153, 157, 148, 145, 149, 151, 137, 151, 157, 147, 144, 140, 142, 135, 150, 147, 141, 147, 127, 138, 129, 141, 140, 137, 139, 151, 139, 146, 147, 140, 141, 154, 149, 157, 160, 160, 152, 153, 146, 139, 153, 149, 151, 151, 125, 132, 137, 135, 127, 127, 130, 115, 138, 142, 141, 153, 154, 159, 146, 151, 154, 161, 151, 150, 157, 147, 149, 146, 161, 160, 151, 141, 144, 151, 143, 149, 148, 146, 152, 145, 151, 143, 144, 150, 139, 138, 147, 140, 146, 153, 143, 149, 150, 151, 155, 140, 129, 151, 155, 157, 153, 147, 153, 152, 153, 154, 141, 136, 136, 148, 148, 152, 138, 141, 132, 143, 128, 129, 149, 140, 139, 137, 138, 137, 141, 150, 140, 139, 131, 139, 143, 139, 135, 142, 135, 134, 135, 133, 121, 116, 120, 123, 122, 117, 101, 109, 114, 110, 107, 111, 115, 124, 121, 119, 131, 139, 126, 117, 124, 133, 131, 115, 126, 126, 117, 120, 108, 121, 124, 121, 126, 130, 125, 128, 138, 139, 137, 128, 124, 125, 145, 130, 130, 138, 133, 150, 144, 143, 147, 140, 150, 138, 142, 130, 128, 131, 139, 135, 131, 136, 139, 133, 136, 139, 133, 127, 121, 120, 135, 132, 136, 136, 126, 134, 123, 130, 140, 131, 135, 141, 149, 157, 144, 153, 153, 147, 159, 141, 148, 141, 139, 149, 136, 145, 145, 125, 125, 137, 155, 141, 134, 148, 147, 150, 147, 142, 149, 152, 156, 150, 157, 149, 147, 153, 151, 149, 150, 150, 155, 146, 146, 156, 150, 148, 150, 144, 147, 152, 146, 130, 155, 156, 134, 150, 148, 141, 139, 135, 140, 144, 139, 134, 135, 148, 146, 149, 144, 156, 157, 153, 145, 164, 160, 156, 152, 149, 155, 146, 139, 144, 139, 140, 128, 129, 132, 131, 131, 133, 138, 141, 146, 148, 159, 151, 149, 154, 155, 159, 140, 158, 160, 156, 151, 146, 154, 150, 150, 155, 148, 149, 146, 151, 145, 141, 141, 130, 142, 145, 153, 148, 155, 156, 152, 147, 148, 154, 151, 141, 152, 159, 159, 148, 144, 153, 151, 144, 152, 148, 147, 148, 138, 141, 147, 144, 144, 141, 139, 145, 135, 139, 143, 140, 138, 132, 145, 140, 136, 143, 145, 138, 137, 139, 144, 145, 144, 143, 148, 142, 128, 133, 126, 132, 125, 125, 131, 127, 129, 118, 121, 125, 117, 105, 107, 118, 109, 112, 116, 117, 126, 118, 124, 133, 131, 125, 119, 132, 133, 100, 115, 116, 119, 132, 124, 120, 123, 124, 125, 122, 120, 128, 140, 142, 133, 134, 129, 120, 135, 134, 134, 136, 126, 128, 134, 146, 137, 144, 133, 138, 135, 131, 127, 124, 131, 132, 133, 132, 143, 130, 135, 131, 129, 136, 142, 137, 128, 132, 132, 118, 132, 135, 115, 140, 160, 140, 137, 144, 147, 146, 153, 147, 141, 137, 158, 144, 147, 149, 147, 141, 141, 146, 146, 149, 137, 155, 148, 147, 142, 138, 151, 142, 145, 154, 154, 152, 148, 156, 138, 150, 144, 158, 150, 147, 150, 147, 144, 147, 141, 141, 152, 146, 164, 145, 136, 143, 253, 148, 152, 147, 148, 148, 142, 148, 139, 139, 141, 140, 136, 140, 153, 138, 149, 147, 155, 148, 156, 154, 146, 159, 160, 157, 158, 152, 147, 138, 147, 151, 145, 134, 130, 139, 123, 122, 137, 139, 136, 152, 146, 147, 153, 153, 161, 156, 157, 157, 154, 149, 154, 160, 148, 157, 163, 153, 159, 160, 137, 149, 151, 141, 135, 130, 151, 129, 155, 138, 146, 148, 149, 149, 157, 156, 143, 146, 155, 149, 142, 149, 154, 148, 151, 151, 149, 155, 144, 150, 144, 145, 137, 152, 138, 147, 151, 144, 145, 137, 139, 133, 138, 141, 138, 139, 145, 135, 117, 140, 142, 130, 132, 135, 146, 149, 147, 152, 150, 151, 147, 134, 134, 127, 125, 124, 120, 123, 123, 126, 128, 133, 133, 112, 110, 109, 106, 105, 111, 113, 119, 124, 129, 134, 133, 124, 124, 132, 122, 115, 118, 112, 120, 127, 110, 129, 125, 114, 117, 123, 125, 131, 129, 128, 133, 132, 138, 127, 137, 124, 109, 157, 135, 134, 139, 144, 137, 140, 143, 141, 129, 143, 118, 130, 134, 134, 136, 131, 132, 134, 143, 131, 136, 138, 141, 131, 135, 130, 126, 145, 132, 140, 113, 134, 135, 125, 144, 145, 147, 140, 137, 142, 147, 149, 147, 144, 147, 140, 148, 143, 145, 141, 155, 150, 152, 157, 118, 151, 137, 146, 144, 150, 147, 148, 157, 154, 151, 151, 143, 152, 153, 152, 159, 149, 142, 146, 135, 146, 142, 151, 150, 132, 152, 146, 140, 158, 147, 144, 146, 152, 150, 145, 150, 146, 152, 142, 140, 144, 133, 147, 164, 160, 149, 149, 149, 149, 155, 151, 154, 165, 162, 157, 153, 150, 149, 149, 135, 141, 143, 130, 129, 132, 124, 128, 141, 141, 144, 151, 157, 148, 152, 154, 148, 147, 160, 158, 155, 154, 157, 163, 161, 150, 150, 152, 151, 157, 155, 151, 149, 150, 126, 140, 158, 163, 152, 149, 154, 156, 153, 145, 155, 156, 149, 150, 149, 149, 143, 143, 145, 147, 148, 156, 162, 155, 160, 152, 146, 151, 148, 148, 151, 146, 150, 146, 149, 140, 134, 145, 135, 141, 137, 147, 140, 144, 134, 133, 138, 126, 130, 143, 149, 154, 152, 151, 149, 142, 151, 140, 134, 127, 117, 121, 136, 141, 154, 153, 168, 175, 179, 161, 142, 114, 108, 98, 102, 108, 111, 138, 129, 131, 114, 124, 129, 126, 117, 110, 103, 111, 127, 124, 114, 116, 113, 114, 117, 126, 132, 128, 131, 126, 129, 117, 139, 138, 137, 138, 118, 125, 141, 139, 135, 132, 149, 136, 142, 135, 135, 134, 132, 145, 132, 139, 138, 148, 134, 139, 140, 144, 134, 138, 139, 156, 134, 122, 132, 138, 132, 143, 136, 142, 134, 141, 145, 150, 142, 140, 136, 151, 140, 150, 152, 149, 143, 137, 148, 140, 144, 138, 150, 152, 138, 130, 151, 169, 142, 145, 146, 154, 144, 151, 155, 151, 150, 156, 157, 157, 147, 157, 158, 148, 158, 148, 144, 139, 148, 152, 149, 142, 147, 149, 149, 150, 151, 140, 155, 139, 149, 151, 157, 147, 141, 142, 150, 146, 134, 152, 169, 167, 160, 145, 148, 158, 152, 161, 147, 160, 153, 152, 149, 156, 149, 149, 139, 145, 135, 131, 128, 128, 132, 137, 141, 137, 134, 149, 148, 157, 151, 145, 155, 138, 147, 164, 158, 161, 157, 155, 158, 160, 164, 155, 153, 150, 159, 160, 158, 146, 109, 133, 166, 191, 189, 152, 149, 145, 149, 149, 149, 157, 155, 148, 156, 139, 134, 146, 134, 167, 146, 157, 159, 152, 161, 159, 162, 148, 150, 156, 151, 148, 138, 147, 154, 144, 142, 142, 130, 147, 139, 148, 143, 146, 144, 134, 145, 133, 133, 138, 148, 159, 161, 162, 156, 152, 145, 137, 128, 126, 121, 125, 132, 142, 159, 163, 181, 197, 211, 204, 204, 168, 125, 109, 105, 103, 92, 133, 126, 115, 120, 115, 130, 91, 104, 119, 119, 130, 127, 121, 123, 117, 125, 117, 122, 113, 119, 128, 128, 130, 140, 141, 136, 139, 128, 134, 136, 123, 142, 144, 141, 134, 129, 144, 131, 140, 135, 140, 145, 138, 146, 146, 135, 144, 150, 125, 141, 146, 140, 139, 129, 151, 130, 138, 131, 118, 127, 121, 130, 154, 136, 138, 128, 138, 142, 129, 148, 140, 154, 142, 146, 148, 149, 152, 144, 147, 146, 144, 149, 145, 156, 136, 141, 156, 156, 152, 157, 153, 140, 154, 153, 146, 151, 145, 155, 152, 149, 151, 154, 142, 156, 154, 151, 148, 147, 156, 152, 149, 148, 141, 146, 142, 155, 145, 149, 126, 145, 151, 159, 144, 149, 157, 144, 127, 116, 142, 174, 158, 151, 142, 148, 153, 148, 146, 150, 152, 149, 147, 159, 159, 158, 155, 156, 138, 129, 119, 133, 125, 131, 139, 138, 137, 140, 143, 155, 153, 163, 135, 145, 153, 157, 150, 161, 167, 158, 152, 162, 161, 158, 160, 153, 157, 151, 150, 154, 136, 102, 137, 171, 189, 196, 136, 148, 157, 143, 147, 152, 149, 152, 146, 147, 143, 143, 149, 145, 147, 150, 158, 149, 149, 153, 155, 150, 150, 149, 138, 153, 150, 139, 140, 153, 146, 140, 135, 150, 148, 134, 149, 144, 152, 151, 142, 145, 151, 153, 140, 152, 155, 164, 164, 157, 156, 136, 120, 107, 115, 114, 114, 126, 139, 154, 170, 178, 189, 206, 222, 231, 218, 196, 146, 116, 114, 103, 105, 120, 109, 105, 97, 147, 108, 118, 125, 124, 126, 127, 126, 118, 121, 113, 115, 120, 119, 123, 122, 139, 130, 135, 146, 147, 140, 132, 141, 130, 133, 134, 149, 143, 136, 138, 119, 125, 127, 145, 142, 143, 137, 139, 136, 136, 144, 129, 131, 141, 136, 128, 130, 131, 143, 150, 142, 125, 128, 138, 137, 132, 141, 123, 132, 135, 133, 142, 137, 153, 136, 141, 146, 143, 144, 144, 145, 143, 143, 132, 149, 147, 145, 150, 155, 152, 147, 148, 152, 152, 144, 144, 142, 164, 147, 144, 145, 143, 155, 156, 153, 150, 152, 147, 150, 153, 150, 146, 150, 151, 158, 142, 158, 147, 139, 151, 150, 165, 142, 145, 153, 162, 144, 157, 155, 155, 135, 125, 141, 161, 146, 137, 142, 147, 145, 142, 153, 160, 159, 151, 149, 149, 149, 161, 154, 149, 150, 150, 130, 119, 126, 138, 139, 142, 136, 142, 140, 148, 157, 152, 155, 133, 150, 160, 161, 153, 171, 159, 162, 159, 163, 166, 156, 155, 157, 151, 145, 153, 129, 107, 134, 158, 171, 174, 152, 147, 147, 143, 142, 128, 136, 156, 135, 142, 143, 154, 153, 154, 151, 138, 140, 151, 154, 147, 152, 152, 152, 143, 146, 164, 162, 148, 143, 145, 143, 146, 137, 144, 148, 143, 153, 148, 141, 151, 144, 140, 141, 154, 142, 157, 157, 156, 164, 152, 144, 126, 100, 86, 95, 101, 106, 117, 136, 153, 172, 180, 186, 207, 219, 234, 228, 236, 214, 159, 124, 106, 101, 116, 116, 102, 109, 117, 98, 117, 126, 125, 119, 110, 128, 120, 120, 125, 118, 123, 121, 124, 120, 154, 134, 127, 122, 150, 131, 159, 127, 152, 157, 137, 135, 147, 147, 139, 142, 142, 137, 159, 148, 137, 136, 138, 141, 142, 145, 133, 115, 146, 148, 134, 137, 108, 136, 149, 139, 135, 140, 135, 134, 133, 139, 131, 134, 135, 140, 150, 141, 144, 140, 140, 135, 129, 141, 136, 135, 136, 133, 137, 131, 138, 138, 143, 147, 145, 146, 146, 146, 149, 145, 152, 143, 150, 146, 151, 146, 148, 149, 153, 147, 150, 152, 147, 153, 143, 147, 148, 151, 158, 155, 150, 140, 148, 156, 150, 138, 143, 139, 164, 161, 167, 159, 137, 155, 155, 148, 158, 153, 153, 145, 145, 151, 140, 138, 135, 132, 160, 162, 147, 137, 137, 147, 148, 150, 149, 155, 163, 146, 136, 140, 144, 149, 141, 142, 142, 147, 142, 162, 149, 155, 150, 157, 158, 153, 147, 174, 162, 159, 164, 158, 166, 168, 165, 158, 156, 161, 157, 161, 128, 144, 155, 168, 160, 149, 135, 130, 135, 124, 143, 140, 143, 129, 151, 136, 155, 158, 155, 156, 132, 151, 152, 155, 149, 152, 150, 161, 126, 144, 167, 184, 165, 147, 150, 147, 135, 133, 152, 141, 131, 143, 145, 139, 155, 157, 148, 153, 149, 150, 157, 156, 158, 162, 150, 127, 93, 76, 86, 86, 90, 103, 115, 132, 151, 181, 191, 185, 200, 219, 228, 235, 243, 236, 222, 161, 112, 106, 108, 118, 121, 129, 115, 126, 119, 131, 115, 127, 106, 120, 132, 127, 127, 122, 119, 116, 125, 126, 132, 122, 145, 137, 142, 92, 182, 147, 131, 133, 130, 142, 132, 154, 143, 140, 145, 145, 141, 140, 143, 136, 146, 143, 149, 144, 141, 127, 136, 138, 132, 140, 127, 137, 133, 134, 131, 141, 139, 136, 128, 137, 137, 144, 137, 146, 138, 142, 136, 133, 134, 134, 134, 136, 130, 135, 142, 130, 131, 137, 132, 131, 138, 147, 150, 137, 150, 154, 148, 153, 141, 139, 142, 148, 145, 138, 141, 148, 148, 148, 137, 167, 146, 147, 151, 149, 139, 145, 159, 153, 145, 145, 145, 152, 149, 153, 141, 132, 158, 164, 158, 153, 138, 156, 157, 155, 143, 160, 151, 155, 147, 148, 141, 131, 130, 117, 154, 169, 149, 139, 121, 139, 138, 145, 148, 159, 159, 149, 138, 140, 145, 167, 149, 145, 138, 135, 144, 155, 157, 148, 163, 158, 159, 159, 153, 168, 162, 149, 169, 157, 163, 165, 160, 165, 152, 167, 164, 162, 165, 149, 155, 155, 154, 151, 141, 146, 147, 143, 144, 149, 148, 143, 144, 148, 142, 148, 166, 153, 144, 153, 156, 154, 140, 153, 157, 149, 128, 145, 167, 174, 162, 147, 148, 153, 139, 136, 149, 150, 150, 149, 146, 154, 149, 158, 159, 147, 145, 152, 165, 168, 174, 153, 130, 104, 78, 77, 84, 89, 98, 86, 114, 139, 152, 168, 178, 194, 211, 220, 227, 241, 249, 246, 243, 215, 153, 121, 105, 121, 122, 118, 116, 125, 122, 116, 120, 132, 123, 116, 129, 128, 110, 120, 112, 111, 116, 125, 131, 116, 125, 136, 137, 135, 141, 147, 144, 140, 144, 136, 140, 139, 130, 148, 139, 131, 133, 142, 133, 135, 138, 141, 144, 142, 143, 142, 133, 132, 144, 137, 139, 139, 134, 140, 131, 131, 142, 141, 133, 126, 122, 147, 139, 146, 146, 143, 133, 131, 131, 135, 132, 130, 130, 134, 127, 111, 134, 145, 132, 121, 118, 130, 129, 132, 140, 149, 142, 138, 136, 141, 139, 137, 127, 122, 129, 126, 146, 148, 150, 151, 151, 150, 142, 148, 142, 143, 151, 149, 149, 155, 148, 155, 155, 156, 147, 134, 150, 158, 148, 155, 148, 148, 155, 147, 146, 156, 144, 149, 137, 144, 149, 130, 149, 125, 129, 146, 139, 132, 145, 144, 137, 136, 153, 159, 153, 145, 138, 149, 153, 162, 156, 147, 138, 138, 154, 155, 159, 153, 161, 163, 165, 163, 158, 159, 161, 163, 150, 153, 154, 158, 167, 168, 160, 159, 165, 159, 165, 164, 171, 157, 152, 157, 141, 148, 141, 147, 147, 151, 138, 143, 150, 139, 148, 157, 151, 157, 149, 152, 156, 147, 157, 151, 146, 141, 128, 137, 159, 157, 152, 153, 145, 148, 149, 143, 138, 149, 145, 143, 141, 155, 153, 152, 155, 159, 161, 157, 162, 170, 166, 135, 105, 70, 67, 70, 76, 79, 98, 89, 117, 141, 137, 147, 177, 193, 215, 219, 236, 231, 240, 244, 241, 238, 190, 135, 117, 116, 119, 131, 123, 130, 130, 128, 117, 133, 132, 128, 126, 131, 131, 128, 120, 120, 102, 117, 121, 107, 124, 126, 138, 143, 137, 132, 141, 140, 141, 138, 138, 140, 127, 142, 138, 147, 137, 135, 144, 149, 143, 134, 145, 142, 138, 135, 144, 141, 127, 125, 142, 144, 140, 148, 139, 134, 146, 139, 134, 129, 131, 132, 138, 138, 133, 129, 136, 130, 134, 138, 128, 144, 138, 147, 139, 126, 129, 122, 117, 120, 114, 125, 118, 128, 131, 144, 140, 143, 141, 129, 127, 134, 125, 127, 132, 122, 136, 138, 140, 150, 143, 138, 146, 144, 153, 150, 150, 153, 113, 173, 145, 147, 137, 164, 150, 151, 169, 164, 153, 144, 157, 156, 150, 140, 155, 153, 147, 144, 149, 147, 149, 139, 147, 148, 138, 134, 126, 126, 147, 146, 149, 137, 142, 154, 148, 142, 128, 148, 146, 156, 156, 148, 141, 148, 152, 141, 167, 162, 158, 158, 160, 161, 159, 162, 172, 157, 132, 152, 157, 149, 160, 163, 163, 164, 166, 162, 164, 162, 163, 166, 167, 151, 148, 139, 139, 143, 139, 144, 147, 153, 149, 156, 136, 149, 148, 150, 150, 139, 147, 157, 149, 149, 143, 149, 142, 134, 129, 152, 143, 158, 146, 149, 154, 145, 143, 146, 157, 137, 149, 149, 154, 161, 153, 161, 159, 165, 168, 166, 159, 115, 82, 56, 68, 64, 74, 76, 91, 91, 100, 120, 133, 150, 179, 196, 211, 223, 234, 238, 239, 247, 243, 243, 221, 161, 120, 118, 111, 122, 113, 126, 129, 133, 133, 127, 130, 133, 127, 130, 129, 125, 122, 122, 130, 114, 128, 130, 125, 130, 143, 138, 138, 131, 140, 137, 132, 139, 133, 134, 137, 139, 133, 135, 141, 151, 139, 145, 147, 147, 141, 147, 147, 145, 143, 137, 137, 124, 133, 137, 134, 144, 122, 147, 140, 115, 126, 146, 135, 145, 136, 135, 127, 133, 135, 133, 125, 134, 129, 139, 128, 148, 150, 145, 145, 131, 119, 116, 118, 123, 125, 122, 121, 125, 134, 138, 133, 123, 119, 122, 125, 130, 126, 125, 129, 130, 142, 139, 137, 143, 137, 132, 138, 146, 158, 152, 154, 157, 150, 154, 143, 160, 139, 151, 166, 155, 157, 148, 155, 151, 145, 150, 156, 159, 143, 146, 149, 147, 151, 155, 147, 139, 149, 129, 120, 118, 121, 133, 145, 142, 141, 144, 130, 151, 139, 150, 148, 148, 152, 147, 148, 155, 152, 155, 157, 149, 167, 165, 158, 165, 168, 165, 168, 115, 123, 192, 202, 153, 163, 159, 154, 165, 158, 162, 168, 161, 169, 176, 174, 144, 149, 138, 143, 145, 146, 149, 149, 143, 151, 149, 147, 150, 149, 149, 149, 150, 153, 149, 149, 144, 145, 153, 145, 156, 140, 143, 150, 145, 149, 137, 146, 148, 145, 158, 152, 139, 137, 155, 152, 155, 158, 166, 165, 171, 177, 168, 145, 108, 69, 49, 57, 60, 66, 78, 95, 73, 94, 107, 138, 155, 174, 189, 206, 220, 236, 244, 247, 245, 248, 243, 243, 178, 128, 115, 122, 128, 121, 120, 133, 139, 136, 130, 130, 143, 128, 139, 129, 137, 130, 128, 137, 120, 121, 130, 126, 128, 140, 144, 137, 142, 148, 130, 131, 132, 133, 134, 153, 133, 138, 129, 125, 136, 134, 131, 141, 138, 137, 143, 136, 142, 138, 133, 138, 126, 136, 141, 133, 135, 126, 123, 132, 137, 127, 130, 143, 130, 128, 121, 124, 139, 136, 123, 120, 118, 129, 128, 126, 153, 160, 154, 154, 136, 119, 116, 120, 122, 123, 120, 112, 120, 123, 125, 128, 126, 124, 124, 121, 112, 117, 124, 119, 120, 130, 132, 137, 131, 130, 128, 133, 138, 150, 150, 150, 149, 148, 150, 146, 148, 143, 141, 158, 160, 153, 154, 150, 154, 146, 147, 166, 155, 156, 143, 148, 145, 156, 157, 148, 136, 144, 131, 136, 126, 113, 114, 136, 139, 140, 148, 136, 160, 145, 151, 140, 152, 148, 145, 152, 150, 152, 154, 160, 154, 153, 166, 161, 161, 163, 173, 164, 77, 103, 213, 229, 146, 160, 164, 169, 174, 166, 158, 157, 174, 167, 162, 168, 146, 145, 149, 144, 149, 149, 150, 148, 153, 153, 159, 130, 171, 152, 156, 153, 151, 156, 146, 148, 144, 151, 157, 152, 145, 152, 154, 150, 150, 146, 147, 148, 144, 141, 149, 147, 147, 149, 157, 158, 154, 164, 166, 168, 170, 178, 172, 132, 88, 53, 47, 52, 49, 54, 68, 77, 87, 89, 107, 127, 152, 173, 190, 206, 224, 240, 247, 240, 240, 237, 243, 240, 201, 127, 111, 124, 119, 125, 129, 129, 125, 133, 133, 124, 142, 129, 124, 124, 138, 133, 136, 135, 122, 124, 131, 131, 124, 137, 126, 136, 132, 151, 158, 171, 131, 115, 131, 143, 135, 123, 123, 123, 139, 138, 141, 148, 136, 143, 140, 136, 134, 138, 147, 140, 140, 129, 142, 125, 131, 132, 117, 124, 127, 132, 134, 132, 128, 129, 125, 132, 140, 137, 133, 124, 131, 137, 119, 140, 161, 160, 156, 155, 151, 126, 113, 118, 121, 134, 118, 115, 121, 112, 107, 122, 125, 123, 120, 117, 115, 113, 112, 117, 122, 124, 122, 131, 122, 124, 118, 123, 137, 137, 150, 152, 143, 149, 150, 149, 152, 137, 147, 158, 159, 152, 154, 153, 154, 150, 138, 148, 161, 147, 148, 144, 143, 150, 149, 129, 121, 122, 151, 177, 160, 111, 89, 150, 174, 133, 142, 136, 165, 154, 156, 154, 150, 145, 139, 144, 166, 159, 159, 161, 162, 150, 173, 164, 164, 168, 172, 172, 105, 94, 164, 190, 164, 173, 167, 170, 168, 171, 163, 167, 160, 162, 132, 190, 148, 150, 153, 148, 148, 142, 142, 148, 150, 156, 154, 158, 158, 149, 158, 156, 158, 147, 140, 143, 151, 153, 149, 149, 148, 148, 152, 154, 147, 148, 144, 159, 144, 144, 143, 148, 142, 146, 149, 151, 155, 159, 170, 167, 176, 178, 164, 121, 64, 41, 27, 45, 51, 55, 69, 71, 87, 82, 98, 125, 158, 174, 186, 203, 226, 244, 241, 239, 246, 243, 245, 240, 221, 137, 119, 126, 122, 125, 125, 129, 145, 110, 134, 137, 137, 131, 129, 139, 129, 128, 131, 140, 131, 121, 133, 138, 127, 130, 125, 126, 122, 119, 130, 164, 150, 134, 133, 132, 139, 137, 172, 119, 122, 131, 132, 138, 140, 146, 141, 137, 133, 124, 160, 142, 134, 138, 141, 121, 117, 148, 156, 136, 131, 138, 132, 127, 126, 133, 133, 128, 135, 140, 139, 141, 135, 142, 141, 160, 169, 170, 167, 162, 156, 121, 124, 126, 127, 117, 114, 119, 108, 87, 64, 107, 115, 126, 121, 114, 109, 105, 110, 118, 113, 111, 128, 112, 118, 126, 111, 108, 131, 145, 146, 149, 151, 154, 149, 154, 151, 145, 142, 158, 156, 147, 153, 150, 144, 168, 160, 141, 150, 160, 153, 141, 150, 144, 146, 103, 103, 116, 159, 194, 165, 108, 84, 135, 173, 135, 147, 133, 154, 158, 164, 145, 156, 151, 151, 151, 152, 155, 148, 158, 161, 164, 166, 163, 163, 170, 161, 162, 177, 136, 153, 160, 161, 168, 159, 165, 167, 172, 171, 159, 162, 159, 128, 174, 166, 152, 149, 144, 143, 148, 137, 139, 167, 154, 148, 147, 150, 154, 161, 159, 156, 154, 143, 147, 148, 151, 144, 152, 145, 150, 157, 154, 151, 148, 141, 148, 151, 148, 150, 145, 147, 156, 148, 157, 160, 161, 170, 172, 169, 181, 151, 110, 51, 23, 25, 35, 49, 57, 64, 69, 70, 79, 96, 120, 152, 169, 192, 209, 228, 241, 239, 240, 245, 242, 246, 235, 235, 163, 122, 125, 131, 127, 119, 129, 142, 131, 140, 142, 141, 127, 127, 144, 134, 128, 122, 150, 137, 133, 124, 130, 132, 136, 128, 123, 127, 125, 123, 133, 151, 139, 99, 116, 143, 154, 184, 140, 125, 120, 132, 133, 137, 137, 137, 133, 127, 133, 134, 128, 137, 137, 140, 132, 101, 147, 159, 113, 150, 162, 126, 103, 121, 129, 130, 137, 137, 134, 128, 137, 127, 147, 166, 170, 177, 183, 172, 171, 167, 145, 136, 139, 127, 109, 115, 127, 118, 88, 90, 102, 115, 116, 117, 115, 110, 109, 106, 117, 110, 108, 108, 111, 115, 119, 112, 114, 116, 145, 152, 147, 150, 152, 150, 151, 153, 150, 149, 151, 163, 155, 146, 150, 138, 142, 154, 151, 150, 151, 145, 134, 140, 136, 136, 104, 97, 110, 164, 180, 172, 127, 108, 129, 140, 135, 132, 139, 141, 168, 161, 168, 152, 147, 145, 153, 150, 154, 159, 154, 163, 159, 164, 162, 158, 168, 174, 160, 173, 179, 162, 169, 169, 167, 160, 160, 169, 176, 174, 163, 159, 154, 180, 143, 147, 152, 149, 156, 149, 151, 155, 129, 158, 151, 147, 158, 153, 157, 157, 159, 157, 152, 150, 142, 156, 156, 141, 160, 147, 147, 149, 148, 150, 152, 154, 146, 146, 156, 141, 145, 155, 150, 152, 161, 162, 162, 175, 177, 171, 173, 161, 103, 46, 28, 30, 42, 40, 53, 56, 63, 72, 78, 95, 120, 140, 143, 168, 208, 236, 242, 244, 240, 240, 242, 239, 247, 226, 171, 120, 115, 124, 129, 128, 119, 145, 133, 128, 134, 140, 138, 126, 135, 135, 133, 131, 136, 127, 144, 121, 122, 138, 134, 127, 141, 129, 132, 137, 119, 144, 152, 112, 115, 134, 136, 136, 142, 135, 107, 126, 137, 140, 140, 134, 136, 131, 145, 140, 146, 137, 137, 137, 146, 128, 139, 120, 94, 149, 148, 135, 145, 141, 132, 126, 128, 133, 141, 132, 145, 137, 132, 155, 174, 182, 192, 184, 181, 170, 157, 141, 137, 132, 118, 113, 115, 108, 110, 103, 107, 106, 110, 100, 110, 103, 110, 118, 122, 111, 101, 109, 106, 108, 115, 112, 113, 117, 126, 134, 160, 149, 151, 152, 147, 147, 147, 155, 149, 145, 154, 158, 156, 153, 132, 163, 153, 140, 148, 141, 167, 160, 130, 145, 122, 84, 106, 146, 154, 151, 143, 125, 126, 135, 137, 145, 132, 124, 162, 156, 163, 150, 143, 157, 157, 155, 157, 153, 154, 167, 164, 161, 161, 158, 178, 166, 167, 174, 171, 170, 166, 169, 180, 155, 175, 178, 164, 174, 158, 156, 158, 163, 153, 149, 150, 149, 155, 145, 157, 157, 149, 160, 152, 151, 150, 159, 159, 158, 158, 160, 160, 157, 153, 147, 145, 150, 152, 151, 147, 154, 152, 154, 148, 154, 151, 152, 156, 154, 152, 157, 150, 151, 158, 163, 164, 170, 175, 177, 179, 153, 99, 34, 22, 25, 30, 31, 47, 56, 59, 66, 75, 95, 137, 149, 144, 140, 169, 236, 239, 243, 242, 239, 237, 242, 242, 213, 157, 121, 119, 122, 125, 137, 130, 122, 120, 131, 129, 136, 143, 136, 132, 134, 136, 136, 134, 117, 131, 122, 127, 122, 127, 120, 123, 131, 132, 136, 137, 127, 147, 151, 125, 128, 126, 104, 134, 154, 144, 129, 131, 139, 138, 134, 140, 138, 136, 132, 137, 137, 139, 142, 141, 128, 140, 147, 126, 143, 135, 135, 139, 128, 139, 130, 135, 138, 142, 138, 144, 141, 147, 161, 176, 180, 182, 187, 175, 177, 167, 143, 143, 128, 117, 113, 115, 116, 106, 98, 101, 100, 107, 109, 108, 107, 113, 103, 116, 109, 100, 88, 107, 98, 102, 107, 115, 116, 130, 133, 160, 154, 153, 141, 152, 145, 148, 144, 145, 139, 146, 154, 154, 157, 142, 160, 149, 147, 126, 123, 177, 170, 147, 135, 133, 113, 119, 128, 130, 124, 151, 135, 122, 138, 153, 149, 147, 139, 144, 155, 157, 160, 146, 161, 151, 157, 160, 168, 165, 170, 157, 169, 158, 156, 168, 158, 168, 170, 172, 167, 169, 167, 172, 163, 169, 173, 163, 168, 164, 149, 154, 168, 156, 150, 152, 147, 145, 147, 154, 156, 143, 158, 156, 151, 153, 157, 158, 157, 163, 151, 154, 147, 154, 150, 150, 153, 146, 154, 148, 157, 157, 153, 156, 148, 153, 147, 150, 151, 157, 153, 161, 169, 158, 161, 164, 167, 170, 171, 183, 150, 96, 41, 24, 19, 31, 27, 48, 56, 51, 60, 74, 89, 138, 153, 147, 128, 143, 200, 232, 237, 244, 241, 240, 244, 239, 206, 140, 114, 126, 110, 130, 138, 130, 121, 127, 126, 139, 136, 148, 128, 132, 136, 138, 131, 132, 138, 136, 125, 125, 134, 127, 130, 141, 134, 123, 129, 148, 123, 134, 141, 160, 137, 134, 112, 115, 132, 153, 148, 139, 143, 131, 143, 138, 128, 144, 135, 148, 138, 127, 143, 135, 143, 135, 144, 137, 111, 148, 133, 147, 138, 142, 142, 144, 147, 139, 143, 148, 134, 139, 167, 170, 188, 187, 186, 182, 178, 165, 155, 142, 137, 120, 113, 116, 104, 103, 98, 104, 109, 101, 105, 103, 100, 108, 103, 104, 110, 92, 82, 94, 95, 100, 104, 99, 98, 125, 137, 138, 149, 153, 143, 148, 142, 154, 152, 144, 145, 146, 148, 146, 146, 165, 147, 150, 147, 141, 119, 145, 145, 129, 129, 126, 131, 124, 140, 141, 130, 142, 130, 126, 144, 153, 146, 151, 144, 149, 148, 150, 160, 185, 155, 150, 160, 153, 164, 171, 157, 149, 180, 189, 171, 159, 158, 155, 166, 173, 165, 166, 173, 170, 167, 173, 170, 171, 165, 163, 156, 164, 160, 173, 156, 137, 143, 152, 149, 150, 150, 160, 149, 146, 151, 155, 157, 154, 160, 161, 158, 158, 150, 149, 148, 149, 149, 140, 151, 143, 151, 152, 154, 142, 152, 158, 152, 153, 152, 154, 156, 150, 164, 165, 164, 170, 165, 166, 178, 185, 148, 110, 39, 23, 20, 34, 36, 51, 56, 55, 61, 70, 93, 138, 157, 145, 144, 159, 189, 209, 231, 240, 237, 241, 245, 235, 208, 132, 118, 109, 114, 123, 131, 127, 132, 131, 138, 140, 131, 144, 136, 130, 135, 128, 139, 138, 151, 132, 133, 126, 141, 124, 131, 134, 143, 134, 133, 134, 123, 131, 132, 142, 133, 158, 131, 108, 124, 147, 134, 132, 142, 129, 134, 142, 142, 139, 118, 143, 142, 135, 125, 125, 151, 140, 132, 146, 138, 142, 142, 131, 134, 141, 143, 143, 144, 140, 149, 148, 155, 144, 174, 174, 185, 185, 188, 183, 181, 183, 159, 151, 143, 134, 117, 111, 101, 101, 103, 105, 105, 99, 100, 104, 105, 99, 100, 90, 88, 83, 83, 84, 87, 89, 94, 98, 115, 117, 147, 144, 131, 149, 145, 140, 142, 142, 152, 139, 143, 149, 152, 146, 157, 160, 148, 147, 150, 152, 137, 154, 133, 107, 135, 134, 144, 133, 138, 138, 133, 149, 139, 135, 127, 146, 147, 141, 146, 142, 146, 145, 149, 173, 162, 161, 153, 149, 159, 150, 152, 146, 168, 187, 170, 158, 174, 164, 170, 167, 162, 166, 168, 177, 165, 165, 171, 167, 175, 168, 158, 169, 158, 170, 156, 147, 147, 151, 136, 144, 151, 149, 148, 147, 148, 139, 143, 152, 150, 161, 159, 151, 155, 152, 151, 150, 150, 155, 151, 144, 149, 149, 138, 149, 154, 159, 149, 159, 153, 151, 157, 153, 168, 154, 166, 170, 169, 173, 186, 184, 154, 109, 47, 19, 24, 34, 39, 46, 53, 65, 60, 66, 91, 123, 162, 155, 149, 164, 185, 198, 218, 232, 233, 237, 233, 233, 184, 130, 117, 116, 143, 126, 128, 129, 139, 129, 136, 146, 138, 144, 142, 136, 140, 137, 137, 135, 135, 132, 125, 139, 137, 137, 121, 143, 144, 136, 130, 150, 135, 133, 145, 121, 126, 166, 148, 123, 148, 171, 138, 140, 161, 128, 132, 132, 139, 143, 122, 139, 130, 136, 133, 138, 135, 143, 149, 147, 135, 152, 140, 143, 137, 146, 146, 155, 152, 141, 146, 150, 151, 157, 177, 180, 190, 189, 183, 182, 188, 183, 174, 163, 149, 131, 123, 105, 112, 105, 105, 91, 96, 100, 100, 98, 97, 95, 83, 78, 81, 76, 73, 68, 77, 79, 83, 96, 110, 123, 138, 134, 137, 145, 143, 133, 148, 138, 153, 136, 136, 148, 157, 147, 156, 148, 158, 150, 148, 156, 148, 150, 146, 133, 132, 140, 148, 154, 135, 144, 140, 153, 146, 140, 128, 131, 137, 144, 146, 151, 141, 141, 154, 155, 157, 155, 149, 159, 157, 155, 141, 139, 162, 178, 161, 151, 167, 164, 172, 161, 174, 169, 165, 173, 166, 168, 176, 171, 169, 169, 162, 174, 170, 167, 156, 156, 136, 150, 151, 147, 149, 151, 155, 154, 150, 147, 152, 152, 153, 159, 157, 158, 156, 149, 146, 146, 149, 152, 143, 148, 146, 144, 150, 151, 150, 153, 131, 165, 153, 154, 161, 164, 173, 165, 170, 164, 173, 171, 170, 182, 159, 122, 58, 22, 13, 37, 50, 51, 51, 52, 69, 71, 90, 109, 138, 153, 155, 169, 194, 201, 212, 226, 231, 239, 239, 225, 164, 123, 110, 121, 126, 126, 143, 140, 137, 131, 140, 143, 147, 131, 133, 139, 151, 146, 131, 133, 126, 134, 131, 138, 141, 138, 132, 130, 132, 126, 136, 132, 131, 141, 136, 121, 101, 148, 132, 114, 148, 183, 132, 116, 169, 151, 150, 131, 129, 133, 145, 138, 142, 137, 135, 137, 138, 141, 138, 142, 139, 146, 140, 146, 151, 144, 148, 151, 141, 151, 148, 149, 152, 164, 183, 179, 189, 195, 199, 195, 196, 186, 180, 170, 151, 139, 124, 109, 108, 111, 104, 104, 89, 88, 94, 97, 90, 88, 90, 73, 70, 67, 57, 68, 65, 64, 77, 79, 90, 121, 127, 126, 122, 127, 141, 139, 142, 140, 146, 145, 139, 148, 152, 152, 152, 149, 150, 157, 154, 153, 140, 145, 152, 147, 126, 146, 140, 155, 146, 139, 151, 149, 148, 151, 129, 135, 133, 130, 145, 149, 144, 152, 153, 145, 159, 164, 152, 159, 158, 154, 144, 142, 154, 153, 159, 151, 157, 161, 170, 172, 169, 162, 165, 165, 173, 169, 167, 170, 163, 175, 166, 175, 169, 163, 155, 147, 154, 163, 153, 148, 145, 154, 149, 158, 154, 152, 148, 156, 147, 156, 159, 156, 157, 146, 151, 152, 158, 147, 156, 149, 149, 152, 157, 150, 152, 154, 150, 158, 178, 189, 185, 191, 180, 163, 165, 164, 169, 180, 179, 179, 161, 137, 92, 39, 26, 35, 51, 48, 44, 51, 50, 74, 79, 94, 119, 136, 153, 166, 182, 195, 207, 212, 228, 235, 228, 194, 158, 124, 111, 129, 133, 126, 131, 145, 139, 133, 130, 141, 144, 139, 138, 134, 142, 142, 134, 126, 134, 148, 136, 139, 138, 137, 139, 139, 127, 129, 129, 128, 132, 139, 138, 140, 123, 123, 109, 109, 153, 159, 143, 120, 113, 147, 179, 136, 128, 131, 141, 131, 140, 146, 137, 142, 138, 141, 142, 133, 151, 136, 146, 140, 148, 142, 139, 142, 140, 148, 141, 145, 144, 158, 181, 185, 194, 186, 192, 197, 199, 194, 197, 167, 148, 139, 135, 131, 134, 122, 102, 94, 87, 94, 79, 78, 82, 86, 87, 66, 60, 52, 51, 43, 50, 59, 63, 70, 93, 110, 119, 122, 125, 121, 134, 139, 138, 140, 143, 144, 148, 148, 156, 152, 153, 161, 152, 153, 158, 157, 142, 147, 140, 141, 135, 152, 148, 143, 149, 151, 146, 154, 150, 147, 147, 143, 133, 133, 148, 148, 145, 138, 143, 136, 155, 166, 149, 150, 161, 166, 159, 144, 155, 161, 159, 167, 159, 163, 164, 164, 168, 168, 161, 165, 170, 167, 172, 174, 163, 171, 168, 175, 176, 162, 147, 152, 149, 145, 152, 157, 151, 151, 155, 154, 152, 156, 158, 156, 157, 150, 151, 144, 160, 152, 132, 156, 162, 153, 141, 154, 151, 154, 145, 149, 158, 154, 149, 148, 150, 157, 151, 163, 161, 165, 164, 158, 173, 173, 177, 176, 172, 141, 109, 64, 30, 34, 44, 43, 55, 62, 67, 68, 76, 96, 110, 131, 145, 160, 176, 180, 206, 210, 215, 229, 214, 155, 125, 112, 120, 128, 132, 141, 137, 139, 139, 139, 136, 138, 137, 142, 144, 137, 145, 141, 145, 143, 132, 134, 129, 131, 136, 134, 147, 133, 124, 127, 134, 138, 129, 135, 135, 144, 134, 141, 126, 107, 137, 137, 132, 133, 115, 123, 164, 174, 126, 124, 138, 132, 130, 139, 150, 145, 134, 149, 142, 142, 149, 143, 141, 140, 154, 148, 144, 141, 137, 155, 142, 146, 150, 154, 168, 190, 190, 192, 197, 203, 195, 194, 195, 182, 165, 153, 140, 137, 141, 127, 105, 101, 89, 81, 73, 65, 73, 69, 78, 59, 56, 53, 48, 35, 36, 46, 54, 57, 67, 79, 111, 117, 117, 125, 134, 142, 132, 135, 139, 142, 146, 144, 143, 153, 156, 151, 150, 146, 150, 152, 143, 160, 159, 146, 145, 149, 148, 157, 145, 150, 151, 133, 145, 139, 144, 154, 143, 142, 155, 156, 152, 155, 155, 135, 153, 149, 142, 142, 166, 169, 155, 155, 146, 164, 164, 166, 166, 168, 161, 167, 163, 167, 169, 174, 175, 169, 165, 173, 170, 166, 169, 177, 173, 172, 144, 160, 152, 150, 146, 141, 140, 144, 149, 159, 157, 155, 153, 154, 157, 152, 158, 154, 154, 156, 154, 154, 152, 148, 149, 153, 153, 152, 146, 151, 151, 149, 147, 145, 149, 156, 156, 154, 161, 164, 158, 164, 163, 173, 171, 175, 167, 157, 136, 91, 56, 45, 37, 46, 40, 56, 67, 76, 77, 97, 113, 129, 130, 151, 170, 179, 181, 199, 211, 214, 178, 129, 112, 110, 124, 123, 132, 137, 138, 141, 139, 137, 139, 149, 139, 126, 155, 138, 140, 146, 141, 138, 134, 132, 143, 142, 131, 132, 135, 131, 134, 133, 134, 129, 124, 126, 139, 147, 132, 137, 141, 142, 144, 146, 133, 131, 123, 146, 121, 160, 137, 129, 142, 139, 147, 144, 144, 141, 138, 145, 146, 143, 145, 147, 147, 141, 143, 142, 153, 150, 133, 139, 144, 144, 153, 150, 166, 190, 194, 188, 183, 200, 198, 199, 186, 190, 168, 165, 143, 147, 152, 152, 106, 99, 85, 76, 65, 65, 69, 68, 69, 53, 60, 61, 36, 36, 25, 44, 46, 52, 58, 72, 94, 111, 117, 132, 138, 136, 133, 134, 134, 142, 149, 139, 150, 153, 152, 149, 160, 155, 148, 151, 144, 154, 157, 152, 152, 151, 152, 148, 155, 146, 153, 150, 141, 141, 144, 150, 137, 142, 154, 154, 154, 154, 156, 142, 146, 151, 149, 148, 142, 167, 154, 156, 158, 166, 154, 160, 182, 162, 166, 163, 167, 155, 178, 179, 174, 175, 172, 147, 172, 158, 170, 167, 167, 174, 152, 152, 155, 137, 161, 146, 140, 157, 140, 144, 147, 149, 157, 157, 155, 152, 154, 162, 161, 151, 152, 160, 154, 154, 161, 160, 152, 150, 145, 151, 155, 150, 146, 127, 155, 157, 159, 158, 162, 164, 157, 167, 169, 172, 171, 175, 174, 166, 150, 122, 80, 44, 30, 45, 49, 46, 59, 77, 73, 87, 96, 104, 127, 147, 157, 169, 165, 198, 201, 176, 142, 117, 108, 120, 130, 122, 139, 129, 148, 146, 143, 149, 141, 145, 135, 138, 142, 137, 144, 145, 147, 143, 124, 136, 145, 142, 125, 129, 123, 129, 136, 136, 134, 126, 126, 127, 138, 124, 116, 130, 137, 140, 137, 135, 145, 128, 124, 140, 124, 120, 137, 131, 144, 138, 136, 131, 146, 149, 143, 140, 147, 146, 137, 142, 149, 147, 134, 152, 146, 141, 140, 146, 133, 141, 149, 148, 141, 176, 178, 186, 177, 194, 201, 203, 190, 197, 184, 173, 151, 159, 160, 152, 121, 100, 77, 59, 67, 70, 74, 78, 84, 64, 60, 57, 35, 34, 17, 39, 34, 41, 53, 61, 86, 115, 117, 117, 127, 127, 129, 140, 143, 147, 156, 150, 149, 152, 150, 152, 151, 149, 153, 151, 153, 147, 158, 151, 151, 156, 150, 156, 151, 155, 149, 148, 141, 141, 144, 141, 130, 153, 150, 147, 142, 142, 143, 153, 150, 145, 156, 158, 155, 144, 165, 142, 168, 163, 152, 144, 205, 168, 168, 166, 161, 162, 166, 178, 173, 167, 171, 159, 166, 169, 169, 178, 163, 164, 154, 159, 154, 155, 148, 152, 147, 149, 149, 143, 150, 152, 154, 151, 150, 157, 153, 148, 159, 152, 152, 157, 160, 162, 153, 148, 151, 156, 147, 162, 151, 151, 157, 151, 160, 153, 157, 158, 159, 158, 156, 166, 168, 166, 170, 171, 180, 169, 162, 147, 122, 82, 45, 42, 41, 47, 52, 86, 88, 83, 98, 114, 128, 139, 146, 162, 177, 192, 170, 138, 119, 114, 113, 123, 134, 142, 138, 104, 158, 177, 131, 144, 137, 141, 138, 140, 138, 150, 139, 126, 143, 152, 138, 138, 144, 141, 129, 135, 140, 129, 137, 126, 126, 130, 122, 122, 128, 129, 122, 132, 140, 132, 140, 145, 140, 140, 136, 141, 145, 130, 124, 153, 136, 143, 137, 140, 138, 146, 142, 159, 142, 140, 142, 145, 143, 146, 139, 128, 153, 152, 149, 144, 150, 148, 145, 145, 140, 163, 176, 174, 162, 191, 196, 211, 198, 193, 184, 177, 164, 158, 158, 149, 111, 98, 83, 68, 75, 71, 76, 84, 90, 93, 74, 30, 32, 22, 20, 27, 27, 22, 44, 50, 71, 103, 118, 114, 122, 123, 129, 137, 138, 140, 147, 147, 150, 151, 150, 151, 141, 146, 155, 158, 146, 154, 152, 146, 148, 144, 150, 152, 148, 159, 154, 149, 142, 141, 147, 147, 139, 147, 156, 142, 133, 142, 143, 146, 155, 143, 150, 154, 148, 166, 160, 148, 160, 156, 165, 149, 167, 175, 166, 161, 154, 166, 165, 169, 168, 166, 175, 165, 165, 159, 179, 177, 168, 166, 152, 148, 150, 149, 142, 156, 151, 156, 157, 153, 158, 157, 154, 154, 162, 156, 156, 149, 152, 150, 150, 151, 159, 156, 152, 157, 160, 149, 145, 162, 151, 148, 149, 149, 154, 159, 159, 159, 163, 163, 163, 158, 172, 170, 169, 171, 172, 170, 175, 160, 142, 127, 102, 68, 39, 46, 46, 65, 79, 88, 90, 111, 119, 123, 140, 160, 168, 161, 133, 114, 127, 120, 124, 120, 133, 133, 142, 120, 150, 155, 140, 139, 138, 132, 142, 141, 143, 140, 137, 137, 138, 137, 141, 138, 134, 133, 134, 119, 134, 132, 134, 120, 119, 122, 112, 130, 125, 122, 134, 125, 137, 138, 123, 149, 142, 123, 117, 129, 135, 139, 120, 143, 144, 146, 141, 143, 148, 154, 119, 168, 139, 137, 144, 149, 148, 143, 147, 142, 143, 150, 155, 142, 146, 145, 149, 146, 141, 148, 176, 174, 147, 184, 203, 204, 203, 205, 194, 168, 166, 166, 162, 159, 118, 86, 72, 60, 71, 68, 68, 91, 91, 90, 97, 50, 30, 17, 12, 18, 20, 18, 29, 53, 57, 84, 107, 116, 110, 127, 135, 132, 137, 146, 151, 149, 154, 156, 150, 143, 160, 152, 154, 155, 157, 158, 154, 150, 148, 139, 156, 155, 148, 149, 169, 146, 138, 146, 145, 146, 150, 151, 142, 155, 141, 134, 140, 141, 152, 150, 151, 150, 141, 167, 152, 144, 148, 162, 158, 171, 163, 162, 172, 161, 160, 164, 159, 166, 173, 165, 166, 166, 169, 153, 171, 174, 169, 167, 149, 152, 146, 157, 156, 145, 155, 141, 147, 135, 161, 157, 154, 149, 160, 153, 152, 158, 151, 146, 163, 162, 166, 153, 157, 151, 165, 162, 147, 147, 151, 157, 152, 143, 150, 154, 160, 161, 163, 158, 165, 165, 161, 170, 169, 168, 166, 166, 175, 175, 162, 146, 149, 135, 101, 65, 71, 76, 75, 88, 101, 111, 124, 119, 145, 157, 141, 127, 115, 105, 128, 133, 121, 114, 144, 107, 141, 170, 167, 128, 136, 136, 135, 138, 140, 155, 144, 146, 141, 137, 140, 143, 141, 141, 142, 142, 140, 117, 131, 131, 140, 132, 126, 133, 132, 139, 125, 126, 145, 127, 136, 140, 123, 135, 140, 143, 136, 134, 134, 132, 137, 125, 118, 156, 143, 136, 144, 140, 129, 154, 154, 138, 135, 141, 145, 143, 148, 126, 162, 140, 144, 151, 151, 142, 136, 140, 140, 129, 164, 179, 190, 198, 198, 216, 199, 194, 203, 189, 167, 153, 161, 152, 110, 80, 76, 63, 66, 66, 83, 94, 113, 121, 107, 66, 37, 15, 9, 7, 9, 5, 16, 37, 57, 68, 95, 112, 112, 122, 130, 130, 140, 142, 150, 153, 151, 153, 153, 128, 145, 153, 148, 147, 156, 149, 156, 160, 154, 146, 153, 161, 151, 134, 152, 158, 149, 140, 143, 150, 138, 145, 140, 142, 141, 133, 141, 140, 145, 146, 152, 140, 144, 153, 144, 140, 147, 160, 147, 168, 165, 162, 159, 170, 165, 159, 161, 161, 170, 170, 161, 184, 174, 164, 177, 171, 168, 171, 150, 150, 148, 148, 152, 155, 151, 149, 161, 153, 158, 163, 162, 153, 168, 156, 160, 163, 149, 161, 158, 150, 152, 154, 159, 144, 156, 163, 146, 155, 155, 159, 158, 140, 136, 153, 150, 160, 163, 158, 159, 164, 166, 172, 164, 158, 167, 169, 173, 175, 169, 163, 169, 169, 162, 128, 114, 107, 100, 101, 112, 123, 128, 123, 141, 142, 133, 120, 123, 116, 130, 128, 128, 131, 153, 104, 126, 147, 149, 140, 142, 146, 121, 133, 140, 140, 145, 141, 142, 141, 142, 152, 135, 140, 142, 139, 136, 131, 129, 132, 130, 126, 132, 138, 132, 140, 134, 129, 117, 133, 134, 134, 131, 130, 139, 141, 133, 135, 131, 138, 146, 134, 119, 135, 133, 153, 141, 143, 131, 141, 136, 136, 144, 142, 142, 145, 143, 139, 147, 143, 147, 140, 148, 144, 138, 143, 137, 140, 172, 180, 189, 198, 211, 209, 193, 196, 206, 176, 180, 167, 153, 142, 114, 98, 86, 70, 65, 69, 82, 104, 125, 126, 95, 37, 12, 13, 18, 25, 7, 4, 16, 24, 49, 63, 87, 108, 114, 125, 134, 133, 139, 144, 144, 149, 145, 165, 155, 130, 157, 161, 148, 149, 154, 154, 157, 155, 158, 153, 151, 159, 159, 143, 145, 148, 157, 157, 140, 152, 141, 143, 146, 145, 143, 141, 138, 146, 153, 153, 151, 147, 136, 153, 157, 153, 158, 156, 149, 160, 170, 157, 162, 152, 163, 156, 158, 154, 168, 171, 169, 177, 170, 167, 177, 167, 177, 168, 150, 151, 145, 146, 157, 156, 155, 149, 154, 158, 150, 161, 160, 158, 159, 139, 159, 170, 151, 158, 168, 154, 152, 157, 155, 148, 147, 150, 148, 151, 159, 153, 154, 154, 149, 161, 164, 159, 162, 160, 159, 158, 158, 162, 157, 157, 159, 164, 166, 170, 168, 164, 166, 171, 169, 160, 154, 150, 138, 133, 138, 143, 142, 144, 135, 136, 135, 128, 131, 127, 127, 142, 136, 131, 149, 142, 115, 139, 134, 141, 142, 145, 136, 147, 144, 139, 138, 120, 133, 146, 142, 151, 144, 137, 137, 135, 130, 144, 139, 140, 131, 131, 136, 127, 137, 133, 138, 132, 136, 131, 117, 133, 136, 132, 133, 137, 137, 130, 139, 140, 139, 132, 138, 128, 149, 138, 140, 151, 146, 137, 150, 145, 142, 148, 136, 135, 136, 134, 134, 135, 149, 148, 137, 151, 149, 142, 141, 144, 181, 188, 191, 204, 208, 217, 196, 193, 198, 197, 172, 170, 156, 146, 120, 101, 79, 64, 62, 70, 84, 99, 115, 118, 81, 11, 0, 2, 16, 46, 44, 7, 13, 20, 45, 64, 82, 111, 127, 134, 130, 141, 144, 148, 149, 152, 148, 157, 153, 143, 160, 159, 148, 147, 157, 154, 150, 152, 152, 154, 151, 150, 153, 156, 152, 152, 133, 160, 146, 143, 142, 147, 144, 149, 144, 149, 141, 146, 149, 145, 153, 138, 136, 151, 140, 151, 154, 164, 148, 161, 152, 159, 157, 154, 166, 154, 150, 151, 173, 163, 166, 171, 164, 166, 180, 178, 174, 175, 155, 148, 146, 151, 158, 149, 154, 146, 155, 156, 156, 158, 158, 158, 162, 154, 166, 159, 159, 156, 160, 156, 162, 149, 149, 145, 150, 137, 138, 153, 153, 154, 162, 158, 152, 156, 156, 163, 163, 161, 168, 163, 160, 160, 157, 149, 159, 158, 160, 173, 176, 165, 171, 168, 163, 159, 163, 159, 158, 151, 148, 141, 145, 145, 147, 141, 144, 134, 129, 130, 142, 144, 138, 136, 148, 148, 150, 146, 139, 142, 127, 135, 129, 150, 136, 134, 137, 130, 138, 142, 140, 143, 146, 134, 140, 141, 137, 139, 139, 130, 138, 133, 131, 144, 139, 140, 132, 125, 126, 133, 133, 132, 142, 138, 140, 140, 139, 138, 132, 136, 140, 131, 127, 119, 150, 146, 141, 140, 133, 149, 145, 140, 131, 158, 138, 144, 146, 134, 144, 152, 148, 147, 154, 133, 136, 138, 134, 153, 186, 184, 196, 197, 210, 210, 204, 198, 195, 182, 177, 180, 157, 145, 131, 109, 91, 73, 67, 69, 64, 87, 100, 102, 69, 10, 2, 0, 1, 54, 82, 18, 19, 17, 37, 63, 80, 114, 123, 124, 131, 128, 147, 148, 146, 151, 153, 152, 142, 152, 154, 160, 160, 156, 156, 159, 148, 160, 157, 152, 154, 143, 159, 150, 154, 156, 146, 155, 153, 145, 141, 151, 141, 141, 156, 141, 144, 148, 147, 149, 144, 144, 109, 149, 159, 155, 156, 157, 143, 148, 159, 153, 159, 155, 160, 164, 160, 165, 153, 169, 157, 166, 167, 164, 178, 194, 156, 178, 157, 152, 157, 148, 156, 149, 155, 141, 168, 155, 166, 154, 156, 156, 163, 157, 153, 158, 161, 157, 155, 151, 164, 157, 161, 152, 154, 157, 141, 153, 157, 153, 153, 149, 156, 157, 164, 153, 153, 157, 160, 160, 168, 158, 152, 155, 162, 160, 155, 169, 171, 167, 164, 165, 168, 167, 168, 165, 155, 159, 151, 151, 150, 153, 143, 150, 148, 145, 139, 137, 136, 145, 146, 144, 134, 142, 149, 127, 123, 168, 162, 129, 131, 145, 141, 143, 135, 139, 140, 145, 139, 136, 139, 140, 135, 139, 137, 131, 135, 124, 128, 133, 138, 139, 132, 126, 143, 141, 145, 129, 129, 131, 141, 136, 136, 143, 137, 139, 137, 139, 138, 135, 137, 129, 129, 139, 142, 136, 143, 146, 134, 154, 118, 136, 144, 141, 127, 172, 147, 143, 131, 169, 142, 138, 139, 145, 147, 155, 178, 194, 196, 194, 206, 207, 206, 199, 187, 184, 175, 179, 167, 148, 146, 113, 101, 82, 69, 73, 61, 75, 92, 84, 68, 9, 1, 0, 1, 25, 80, 15, 2, 13, 39, 61, 74, 103, 116, 131, 129, 133, 133, 143, 144, 153, 147, 150, 137, 172, 149, 162, 156, 156, 145, 156, 154, 154, 156, 148, 150, 149, 154, 150, 154, 160, 141, 140, 159, 153, 146, 156, 142, 138, 146, 150, 142, 146, 141, 148, 147, 151, 149, 148, 160, 159, 144, 160, 161, 165, 161, 156, 156, 158, 163, 157, 175, 166, 161, 172, 160, 147, 156, 171, 162, 188, 167, 168, 165, 143, 157, 150, 152, 146, 154, 152, 156, 163, 160, 153, 155, 160, 160, 163, 161, 167, 159, 157, 155, 149, 163, 156, 158, 152, 158, 163, 149, 149, 159, 155, 157, 149, 146, 153, 154, 156, 158, 159, 166, 164, 167, 158, 158, 158, 164, 166, 158, 164, 165, 164, 165, 148, 160, 162, 160, 165, 165, 162, 156, 143, 148, 151, 147, 142, 150, 145, 149, 152, 143, 142, 147, 153, 143, 144, 147, 132, 106, 140, 163, 160, 148, 136, 143, 147, 134, 128, 131, 147, 139, 140, 137, 139, 139, 134, 143, 145, 132, 96, 129, 138, 135, 133, 132, 141, 128, 138, 146, 133, 130, 141, 138, 135, 135, 144, 147, 155, 146, 131, 139, 136, 137, 141, 131, 144, 140, 146, 133, 133, 138, 141, 146, 143, 145, 144, 104, 159, 142, 149, 158, 141, 138, 140, 145, 145, 152, 160, 179, 184, 203, 207, 207, 198, 206, 206, 189, 189, 180, 181, 172, 158, 145, 131, 113, 96, 76, 68, 75, 67, 73, 85, 74, 10, 0, 0, 0, 16, 33, 3, 6, 22, 40, 56, 76, 100, 114, 127, 122, 132, 138, 141, 138, 146, 156, 156, 139, 155, 147, 158, 161, 152, 161, 157, 154, 155, 158, 155, 148, 153, 145, 152, 159, 157, 132, 148, 170, 151, 143, 148, 153, 146, 153, 141, 155, 140, 144, 144, 146, 149, 146, 158, 149, 165, 153, 157, 149, 160, 167, 162, 157, 160, 165, 160, 175, 162, 160, 163, 174, 161, 139, 160, 183, 187, 170, 158, 155, 155, 155, 157, 155, 153, 158, 157, 157, 164, 161, 170, 157, 161, 158, 159, 143, 157, 158, 158, 154, 157, 163, 160, 158, 158, 162, 159, 155, 152, 153, 152, 160, 157, 155, 154, 148, 153, 150, 161, 155, 156, 158, 156, 157, 153, 155, 162, 160, 163, 168, 164, 162, 150, 161, 153, 159, 157, 164, 161, 153, 150, 147, 152, 149, 145, 152, 145, 148, 149, 139, 148, 147, 149, 151, 149, 155, 148, 125, 126, 137, 135, 143, 138, 137, 143, 143, 132, 123, 130, 134, 139, 136, 138, 134, 137, 142, 141, 145, 136, 135, 138, 137, 137, 131, 137, 133, 124, 131, 135, 130, 135, 135, 140, 138, 132, 138, 134, 144, 130, 144, 136, 140, 138, 127, 143, 129, 144, 143, 135, 125, 135, 153, 149, 140, 151, 141, 141, 135, 131, 143, 143, 148, 143, 146, 148, 145, 152, 185, 183, 199, 205, 206, 204, 206, 214, 195, 190, 193, 191, 173, 162, 165, 144, 128, 110, 86, 75, 75, 71, 81, 76, 58, 26, 5, 0, 3, 7, 6, 2, 10, 22, 42, 55, 69, 99, 102, 124, 122, 134, 135, 136, 143, 143, 145, 156, 152, 150, 156, 156, 158, 155, 159, 148, 153, 152, 153, 157, 151, 150, 149, 153, 161, 154, 134, 137, 159, 164, 158, 141, 148, 144, 145, 139, 146, 153, 144, 140, 148, 147, 155, 154, 151, 151, 144, 153, 156, 153, 164, 157, 163, 162, 162, 164, 165, 170, 156, 161, 173, 168, 130, 156, 165, 159, 165, 155, 149, 144, 149, 156, 151, 154, 163, 148, 157, 159, 157, 163, 156, 158, 157, 166, 157, 150, 158, 159, 156, 150, 164, 160, 156, 151, 157, 165, 153, 156, 155, 158, 158, 147, 150, 155, 149, 155, 154, 151, 153, 160, 159, 164, 154, 147, 166, 159, 158, 160, 160, 160, 161, 156, 154, 152, 160, 156, 157, 157, 149, 152, 149, 145, 155, 145, 150, 152, 152, 148, 148, 148, 149, 149, 153, 152, 149, 137, 149, 146, 138, 140, 146, 138, 146, 136, 142, 139, 137, 133, 140, 143, 139, 136, 135, 137, 138, 141, 145, 138, 142, 145, 141, 138, 136, 138, 129, 132, 126, 105, 101, 129, 134, 140, 120, 126, 126, 151, 125, 139, 140, 141, 130, 122, 142, 139, 134, 137, 139, 138, 133, 144, 145, 141, 139, 146, 136, 139, 150, 147, 142, 141, 150, 141, 136, 146, 148, 147, 177, 184, 199, 205, 209, 207, 203, 211, 200, 198, 198, 192, 182, 176, 166, 143, 133, 114, 104, 88, 79, 77, 80, 63, 52, 40, 42, 12, 12, 11, 6, 10, 11, 30, 33, 55, 57, 91, 105, 126, 126, 128, 128, 132, 138, 148, 148, 147, 147, 144, 157, 163, 154, 160, 158, 151, 153, 153, 158, 153, 161, 162, 158, 157, 154, 151, 152, 140, 132, 165, 167, 156, 149, 138, 152, 144, 150, 146, 148, 147, 149, 141, 147, 135, 158, 143, 145, 148, 153, 147, 174, 166, 156, 152, 156, 130, 159, 167, 167, 156, 158, 168, 145, 159, 161, 151, 165, 168, 160, 147, 151, 154, 155, 153, 162, 154, 157, 161, 161, 161, 156, 160, 162, 166, 156, 137, 158, 157, 150, 155, 164, 155, 150, 152, 152, 155, 154, 148, 148, 152, 152, 151, 142, 151, 159, 146, 150, 154, 154, 154, 156, 157, 151, 148, 157, 157, 162, 158, 153, 162, 158, 164, 156, 160, 154, 143, 151, 152, 178, 152, 155, 156, 149, 146, 149, 149, 149, 149, 151, 151, 156, 157, 153, 151, 147, 139, 145, 151, 153, 140, 141, 131, 147, 131, 142, 140, 141, 140, 139, 138, 127, 125, 140, 140, 138, 132, 147, 142, 138, 138, 143, 139, 131, 138, 132, 144, 135, 128, 121, 132, 136, 141, 136, 133, 135, 138, 134, 139, 137, 150, 133, 129, 139, 121, 123, 118, 137, 133, 139, 136, 110, 179, 144, 144, 140, 135, 143, 149, 147, 147, 143, 142, 145, 139, 140, 138, 152, 190, 194, 206, 215, 211, 206, 206, 206, 198, 195, 190, 193, 184, 168, 147, 137, 119, 100, 94, 79, 82, 61, 56, 63, 56, 56, 32, 24, 20, 13, 22, 25, 42, 38, 52, 69, 86, 99, 118, 127, 127, 132, 116, 147, 142, 148, 150, 155, 154, 155, 152, 152, 152, 185, 157, 149, 150, 155, 163, 156, 162, 157, 151, 155, 150, 156, 147, 140, 157, 143, 163, 145, 150, 157, 155, 140, 151, 147, 150, 149, 146, 156, 130, 159, 166, 161, 152, 178, 153, 155, 148, 159, 158, 160, 154, 155, 168, 162, 162, 156, 161, 163, 165, 163, 163, 165, 164, 164, 156, 156, 149, 149, 155, 152, 156, 159, 164, 159, 165, 161, 155, 155, 156, 164, 158, 152, 149, 151, 154, 157, 160, 151, 159, 155, 163, 161, 152, 150, 156, 152, 147, 145, 159, 155, 155, 154, 158, 154, 152, 162, 158, 158, 155, 149, 157, 160, 163, 159, 158, 157, 164, 169, 159, 160, 155, 115, 127, 168, 159, 152, 152, 148, 147, 132, 144, 153, 150, 148, 151, 152, 149, 159, 152, 149, 149, 146, 145, 148, 155, 140, 121, 121, 136, 141, 141, 135, 130, 131, 123, 122, 130, 136, 137, 133, 131, 139, 136, 133, 138, 136, 127, 129, 130, 129, 128, 137, 132, 135, 128, 135, 137, 138, 138, 132, 130, 133, 138, 139, 142, 131, 133, 142, 125, 128, 132, 137, 140, 144, 139, 121, 138, 142, 130, 149, 143, 141, 150, 153, 135, 152, 145, 143, 135, 142, 143, 135, 160, 178, 203, 215, 212, 220, 209, 211, 205, 203, 200, 192, 183, 174, 154, 135, 122, 98, 84, 81, 75, 68, 60, 59, 57, 60, 47, 35, 27, 19, 32, 37, 40, 47, 60, 71, 83, 94, 112, 121, 133, 131, 134, 139, 140, 142, 143, 153, 149, 143, 139, 159, 149, 163, 153, 146, 153, 160, 155, 156, 155, 164, 151, 150, 157, 153, 150, 149, 156, 149, 157, 164, 155, 157, 151, 154, 143, 137, 151, 151, 145, 151, 151, 147, 168, 153, 137, 201, 180, 148, 157, 153, 155, 152, 163, 156, 161, 163, 172, 161, 165, 157, 165, 168, 170, 172, 174, 156, 153, 157, 156, 158, 155, 156, 158, 158, 166, 159, 166, 161, 158, 151, 158, 157, 161, 156, 148, 159, 157, 159, 158, 155, 159, 155, 158, 157, 157, 152, 152, 154, 151, 154, 153, 154, 153, 157, 159, 157, 145, 152, 157, 157, 155, 159, 158, 156, 155, 152, 157, 151, 159, 158, 160, 154, 151, 169, 136, 140, 144, 159, 157, 147, 143, 141, 144, 148, 152, 151, 157, 145, 153, 148, 160, 147, 144, 143, 152, 143, 145, 145, 136, 122, 144, 147, 132, 132, 125, 99, 102, 115, 134, 135, 134, 141, 134, 141, 147, 135, 136, 135, 128, 147, 145, 131, 117, 130, 134, 132, 130, 133, 132, 134, 144, 131, 140, 138, 138, 135, 140, 131, 137, 138, 137, 122, 120, 152, 144, 141, 142, 139, 159, 150, 139, 148, 137, 143, 141, 145, 140, 143, 146, 139, 141, 132, 132, 126, 151, 167, 188, 219, 214, 215, 218, 216, 211, 205, 199, 202, 187, 170, 164, 143, 124, 99, 84, 67, 68, 61, 55, 60, 61, 63, 51, 46, 35, 38, 41, 43, 39, 49, 59, 70, 81, 91, 104, 113, 133, 127, 128, 111, 163, 137, 162, 146, 148, 150, 147, 155, 152, 150, 144, 147, 154, 153, 158, 146, 144, 168, 149, 153, 152, 135, 155, 157, 158, 156, 151, 147, 160, 154, 148, 139, 137, 133, 136, 156, 149, 148, 158, 147, 159, 142, 118, 182, 192, 148, 147, 153, 161, 157, 166, 150, 157, 166, 168, 158, 163, 164, 170, 168, 173, 159, 174, 144, 156, 162, 153, 151, 158, 162, 157, 156, 162, 163, 155, 155, 161, 165, 160, 157, 160, 155, 155, 160, 157, 157, 159, 161, 154, 144, 150, 155, 148, 153, 158, 151, 148, 155, 158, 158, 156, 149, 151, 157, 151, 149, 153, 152, 151, 156, 156, 157, 145, 142, 151, 145, 149, 158, 155, 147, 145, 157, 144, 151, 140, 148, 149, 153, 147, 150, 151, 145, 157, 151, 152, 157, 152, 145, 150, 167, 148, 151, 148, 149, 141, 140, 142, 128, 148, 142, 129, 132, 123, 92, 89, 123, 125, 129, 141, 143, 136, 127, 146, 150, 140, 139, 126, 141, 137, 133, 133, 127, 134, 139, 128, 132, 137, 130, 142, 140, 136, 161, 125, 127, 140, 129, 129, 128, 135, 130, 115, 128, 133, 140, 137, 139, 140, 143, 130, 158, 144, 144, 136, 145, 149, 145, 139, 124, 142, 163, 159, 139, 152, 157, 188, 205, 217, 222, 218, 217, 205, 210, 203, 202, 194, 176, 170, 147, 130, 107, 85, 59, 59, 54, 55, 47, 57, 57, 59, 66, 46, 50, 53, 54, 51, 58, 61, 67, 81, 85, 99, 111, 124, 121, 125, 117, 139, 136, 140, 138, 138, 151, 151, 153, 153, 157, 145, 153, 156, 158, 156, 145, 155, 166, 153, 139, 164, 169, 140, 159, 157, 149, 159, 129, 154, 149, 151, 149, 141, 132, 143, 137, 147, 152, 156, 152, 157, 153, 135, 153, 164, 162, 152, 157, 153, 156, 161, 156, 163, 172, 162, 157, 166, 161, 172, 169, 159, 168, 173, 145, 157, 161, 155, 150, 167, 158, 154, 157, 158, 161, 156, 156, 147, 157, 151, 168, 161, 155, 156, 169, 154, 154, 158, 162, 155, 156, 164, 161, 151, 151, 148, 152, 156, 150, 156, 149, 160, 153, 158, 156, 159, 147, 130, 149, 149, 155, 165, 158, 147, 148, 151, 145, 148, 151, 153, 153, 158, 154, 152, 152, 149, 145, 145, 146, 155, 155, 150, 146, 154, 153, 148, 154, 146, 150, 148, 144, 152, 163, 142, 151, 147, 145, 138, 126, 145, 140, 121, 146, 128, 109, 102, 122, 137, 132, 142, 140, 147, 135, 140, 133, 138, 132, 127, 142, 144, 132, 130, 133, 132, 136, 132, 129, 134, 126, 137, 130, 101, 179, 156, 132, 136, 133, 137, 140, 136, 133, 139, 135, 125, 132, 138, 138, 132, 163, 141, 138, 143, 144, 141, 153, 147, 142, 121, 110, 137, 155, 173, 139, 158, 157, 188, 203, 214, 224, 228, 223, 213, 211, 205, 201, 202, 188, 157, 143, 134, 107, 82, 61, 61, 47, 52, 57, 56, 61, 58, 62, 56, 58, 65, 64, 56, 53, 71, 74, 74, 73, 87, 105, 121, 119, 116, 125, 113, 149, 134, 136, 139, 151, 147, 151, 149, 157, 151, 155, 161, 157, 154, 149, 148, 155, 154, 121, 149, 183, 149, 156, 154, 147, 142, 133, 150, 148, 151, 145, 165, 139, 139, 136, 144, 149, 158, 152, 147, 163, 153, 155, 154, 156, 152, 149, 157, 156, 158, 151, 155, 156, 162, 162, 168, 165, 177, 179, 165, 167, 166, 155, 154, 154, 161, 148, 151, 154, 163, 153, 156, 162, 157, 158, 151, 150, 150, 154, 155, 164, 153, 160, 163, 156, 157, 157, 152, 150, 168, 157, 156, 146, 142, 151, 157, 158, 155, 156, 159, 158, 155, 156, 155, 154, 151, 166, 148, 155, 158, 161, 154, 158, 153, 157, 147, 153, 157, 159, 159, 149, 153, 174, 162, 142, 139, 155, 150, 152, 145, 151, 152, 147, 134, 155, 147, 155, 135, 142, 160, 162, 145, 145, 141, 143, 140, 137, 139, 143, 121, 124, 160, 120, 125, 133, 140, 134, 137, 138, 144, 144, 146, 123, 128, 146, 128, 129, 144, 133, 133, 137, 126, 131, 136, 140, 138, 140, 135, 137, 111, 123, 126, 131, 144, 133, 140, 129, 130, 138, 135, 125, 126, 130, 138, 129, 121, 151, 145, 140, 131, 142, 147, 147, 145, 142, 110, 99, 127, 153, 171, 142, 144, 152, 186, 203, 211, 219, 226, 223, 215, 218, 215, 210, 206, 198, 162, 156, 132, 108, 91, 70, 56, 55, 44, 53, 53, 55, 49, 57, 56, 65, 75, 68, 66, 61, 60, 74, 74, 78, 97, 104, 109, 114, 97, 116, 107, 143, 139, 134, 151, 148, 143, 142, 154, 152, 159, 155, 156, 154, 156, 156, 154, 157, 152, 144, 143, 149, 157, 160, 155, 159, 151, 150, 155, 144, 150, 147, 149, 133, 123, 132, 144, 144, 143, 153, 142, 146, 148, 159, 153, 151, 154, 158, 152, 151, 152, 156, 160, 158, 156, 159, 169, 165, 172, 166, 169, 172, 178, 159, 151, 154, 161, 161, 159, 150, 161, 151, 156, 157, 160, 152, 153, 155, 160, 164, 156, 154, 156, 150, 160, 170, 150, 164, 164, 144, 162, 157, 162, 149, 151, 151, 152, 155, 154, 153, 151, 152, 152, 152, 151, 158, 152, 159, 161, 159, 154, 159, 155, 161, 160, 159, 153, 152, 162, 160, 158, 121, 132, 187, 210, 154, 145, 157, 153, 150, 148, 149, 149, 151, 150, 151, 150, 151, 124, 160, 165, 137, 148, 145, 148, 145, 144, 135, 136, 133, 114, 122, 161, 142, 133, 131, 134, 139, 136, 138, 140, 127, 146, 143, 129, 138, 129, 130, 125, 131, 125, 138, 134, 130, 138, 136, 139, 135, 133, 136, 121, 124, 135, 131, 137, 134, 136, 126, 129, 139, 139, 128, 133, 127, 130, 140, 142, 138, 135, 156, 131, 142, 137, 151, 145, 145, 126, 108, 128, 146, 158, 137, 148, 154, 186, 207, 213, 218, 222, 220, 217, 210, 218, 212, 208, 192, 186, 166, 137, 115, 93, 73, 67, 54, 42, 44, 53, 53, 59, 60, 66, 60, 73, 73, 70, 69, 61, 72, 74, 78, 94, 107, 104, 86, 137, 99, 121, 122, 130, 137, 137, 142, 148, 144, 151, 143, 140, 169, 147, 155, 146, 159, 153, 148, 150, 149, 161, 151, 157, 154, 149, 162, 158, 157, 146, 151, 153, 142, 152, 146, 141, 144, 151, 147, 140, 149, 158, 155, 139, 158, 158, 148, 161, 156, 156, 155, 159, 158, 158, 166, 159, 153, 171, 173, 161, 152, 167, 169, 173, 157, 156, 155, 151, 160, 154, 155, 158, 162, 158, 162, 159, 165, 156, 157, 144, 156, 159, 158, 153, 154, 144, 158, 158, 148, 158, 150, 155, 163, 152, 154, 156, 157, 159, 157, 159, 155, 151, 145, 154, 149, 149, 158, 158, 155, 156, 156, 156, 160, 154, 158, 160, 160, 157, 156, 156, 155, 142, 97, 126, 168, 195, 162, 144, 151, 145, 153, 155, 153, 149, 150, 155, 146, 145, 143, 124, 162, 164, 141, 136, 142, 137, 131, 152, 138, 136, 127, 121, 127, 150, 134, 118, 117, 131, 135, 134, 135, 141, 140, 135, 131, 140, 138, 134, 139, 135, 132, 109, 141, 131, 133, 130, 133, 131, 138, 135, 130, 121, 130, 136, 135, 136, 130, 135, 129, 134, 138, 143, 123, 140, 101, 115, 148, 142, 142, 146, 135, 142, 144, 133, 139, 152, 147, 138, 136, 135, 138, 144, 137, 140, 157, 189, 205, 209, 216, 225, 218, 218, 211, 211, 217, 212, 194, 192, 170, 147, 126, 109, 92, 68, 56, 53, 43, 40, 49, 51, 56, 65, 66, 67, 65, 53, 70, 68, 66, 75, 83, 97, 101, 97, 52, 155, 107, 127, 122, 134, 138, 140, 144, 147, 143, 152, 138, 133, 175, 158, 153, 158, 155, 157, 148, 156, 150, 158, 154, 154, 147, 152, 161, 165, 162, 149, 150, 157, 147, 146, 146, 140, 144, 138, 135, 143, 149, 152, 149, 149, 156, 153, 150, 160, 152, 150, 154, 150, 158, 163, 165, 162, 158, 171, 168, 160, 158, 182, 177, 170, 153, 155, 163, 151, 153, 151, 159, 157, 160, 155, 154, 157, 148, 158, 158, 160, 153, 156, 152, 162, 163, 158, 155, 162, 153, 160, 145, 149, 148, 156, 154, 156, 157, 149, 149, 150, 153, 150, 148, 150, 155, 150, 155, 159, 150, 156, 157, 156, 155, 158, 157, 151, 158, 161, 155, 158, 160, 138, 112, 126, 155, 160, 144, 150, 153, 148, 145, 152, 155, 147, 148, 144, 149, 151, 151, 138, 145, 157, 143, 126, 164, 149, 148, 154, 146, 149, 141, 134, 129, 143, 131, 123, 128, 120, 126, 137, 135, 127, 137, 141, 134, 133, 147, 135, 128, 127, 132, 118, 136, 129, 132, 129, 130, 126, 133, 130, 133, 130, 137, 141, 142, 127, 130, 144, 137, 137, 136, 141, 136, 139, 118, 124, 124, 125, 129, 127, 127, 127, 124, 120, 123, 129, 144, 147, 143, 143, 149, 136, 133, 137, 155, 182, 198, 207, 215, 220, 218, 213, 218, 209, 213, 207, 207, 194, 176, 138, 138, 118, 95, 82, 60, 60, 45, 46, 56, 44, 52, 59, 59, 63, 69, 61, 69, 75, 74, 75, 87, 92, 94, 91, 105, 103, 106, 126, 130, 136, 142, 137, 147, 143, 140, 142, 142, 151, 159, 163, 151, 159, 153, 162, 156, 156, 150, 159, 151, 150, 147, 155, 167, 156, 150, 147, 150, 145, 148, 145, 143, 152, 142, 142, 137, 144, 153, 151, 156, 150, 150, 150, 163, 160, 157, 155, 158, 160, 137, 168, 165, 148, 157, 167, 172, 154, 153, 184, 165, 161, 152, 162, 151, 155, 154, 152, 147, 150, 150, 155, 158, 159, 152, 154, 162, 160, 158, 152, 155, 154, 162, 155, 153, 157, 147, 151, 158, 153, 147, 145, 151, 160, 152, 155, 150, 158, 148, 149, 152, 148, 151, 150, 159, 157, 150, 152, 155, 149, 158, 147, 167, 162, 156, 160, 153, 150, 158, 154, 151, 141, 146, 146, 143, 142, 153, 151, 152, 150, 147, 147, 142, 148, 156, 146, 154, 150, 142, 158, 149, 147, 140, 143, 134, 147, 137, 145, 139, 135, 125, 129, 124, 120, 132, 131, 127, 132, 135, 127, 135, 137, 133, 129, 132, 135, 139, 134, 138, 138, 137, 132, 131, 131, 130, 132, 128, 122, 132, 135, 140, 138, 138, 130, 126, 146, 138, 144, 138, 141, 133, 144, 127, 130, 122, 121, 113, 119, 118, 116, 111, 109, 116, 102, 110, 128, 156, 137, 145, 144, 144, 144, 148, 192, 194, 205, 218, 216, 224, 220, 216, 216, 206, 213, 201, 186, 181, 163, 152, 130, 108, 82, 63, 62, 48, 43, 47, 52, 54, 57, 56, 57, 71, 64, 67, 68, 69, 71, 83, 92, 98, 108, 117, 111, 119, 127, 131, 130, 148, 137, 146, 148, 143, 145, 142, 145, 153, 156, 147, 157, 152, 152, 157, 156, 152, 158, 158, 145, 153, 158, 165, 150, 142, 138, 157, 141, 154, 147, 138, 145, 145, 142, 143, 150, 141, 155, 157, 148, 149, 156, 145, 162, 156, 156, 154, 163, 157, 156, 163, 159, 142, 169, 165, 177, 167, 167, 160, 170, 152, 159, 154, 155, 154, 144, 155, 144, 149, 155, 158, 159, 161, 151, 156, 156, 159, 158, 158, 146, 165, 157, 159, 142, 132, 157, 183, 188, 166, 144, 137, 157, 155, 151, 150, 151, 147, 146, 148, 153, 147, 154, 155, 144, 151, 170, 156, 149, 155, 158, 160, 161, 157, 158, 157, 149, 151, 154, 150, 150, 155, 143, 141, 149, 155, 149, 137, 158, 150, 153, 129, 123, 153, 150, 152, 153, 143, 148, 149, 145, 140, 151, 138, 146, 142, 144, 136, 139, 141, 131, 120, 134, 134, 123, 131, 130, 137, 130, 127, 128, 127, 107, 114, 125, 134, 134, 138, 137, 138, 137, 129, 132, 133, 135, 128, 131, 135, 142, 139, 135, 130, 144, 140, 141, 122, 146, 138, 140, 146, 134, 134, 127, 126, 116, 126, 111, 110, 108, 106, 101, 105, 87, 91, 101, 137, 140, 142, 140, 146, 145, 152, 183, 189, 199, 210, 218, 212, 206, 214, 215, 216, 211, 208, 201, 174, 165, 161, 131, 106, 95, 67, 63, 55, 44, 49, 38, 34, 39, 49, 54, 73, 63, 68, 72, 69, 67, 81, 101, 96, 116, 118, 122, 126, 126, 136, 134, 147, 141, 141, 151, 149, 151, 141, 129, 150, 152, 155, 156, 155, 147, 151, 150, 155, 160, 157, 157, 156, 157, 155, 143, 136, 145, 151, 148, 159, 145, 119, 140, 140, 144, 142, 156, 150, 154, 158, 158, 143, 152, 141, 157, 149, 159, 161, 157, 157, 161, 161, 159, 142, 179, 167, 165, 162, 163, 157, 186, 152, 153, 157, 146, 148, 139, 152, 146, 156, 149, 149, 153, 163, 150, 154, 161, 149, 154, 161, 158, 157, 151, 146, 115, 120, 143, 180, 201, 202, 149, 148, 146, 158, 154, 146, 150, 151, 154, 150, 155, 155, 146, 136, 128, 161, 167, 149, 150, 156, 146, 154, 156, 154, 149, 152, 156, 142, 153, 150, 162, 146, 141, 150, 141, 140, 135, 148, 153, 151, 148, 135, 128, 137, 139, 149, 156, 135, 146, 155, 148, 140, 139, 142, 131, 133, 142, 127, 137, 154, 136, 131, 123, 131, 132, 119, 126, 126, 117, 129, 122, 124, 115, 94, 122, 129, 129, 135, 133, 134, 136, 136, 132, 134, 129, 121, 127, 135, 134, 137, 136, 127, 129, 128, 134, 140, 138, 136, 135, 137, 138, 129, 128, 121, 112, 119, 105, 92, 92, 95, 95, 103, 104, 101, 104, 116, 131, 135, 142, 145, 145, 166, 182, 181, 185, 204, 212, 213, 206, 209, 209, 211, 205, 210, 204, 181, 170, 161, 138, 128, 103, 80, 69, 59, 44, 44, 36, 35, 37, 44, 51, 58, 68, 68, 59, 70, 72, 80, 104, 98, 117, 128, 125, 130, 136, 132, 139, 147, 146, 143, 150, 147, 142, 138, 136, 150, 140, 149, 149, 155, 143, 153, 143, 159, 158, 162, 161, 156, 152, 163, 151, 141, 149, 150, 139, 187, 144, 139, 146, 146, 145, 145, 151, 146, 154, 163, 156, 137, 155, 151, 135, 136, 165, 166, 162, 150, 157, 155, 162, 158, 163, 157, 165, 165, 158, 163, 162, 143, 146, 144, 150, 145, 141, 138, 148, 155, 154, 156, 161, 150, 154, 161, 157, 155, 157, 156, 156, 154, 163, 145, 98, 111, 143, 175, 190, 214, 166, 154, 148, 158, 154, 148, 158, 158, 149, 151, 159, 151, 128, 122, 148, 164, 156, 145, 150, 151, 152, 152, 163, 155, 156, 153, 153, 123, 156, 157, 146, 145, 154, 156, 151, 151, 144, 149, 138, 144, 147, 138, 143, 162, 144, 146, 152, 139, 137, 158, 150, 142, 129, 141, 139, 139, 140, 122, 134, 138, 122, 132, 125, 128, 134, 133, 123, 113, 136, 133, 122, 132, 130, 113, 125, 133, 123, 140, 131, 131, 128, 133, 117, 121, 122, 117, 118, 114, 112, 122, 120, 121, 115, 114, 112, 130, 135, 130, 133, 133, 136, 134, 126, 120, 111, 110, 99, 92, 73, 83, 79, 87, 84, 93, 100, 101, 97, 127, 141, 139, 144, 165, 179, 175, 185, 201, 202, 210, 205, 210, 206, 207, 206, 205, 192, 194, 181, 182, 156, 142, 117, 99, 71, 63, 47, 45, 38, 40, 42, 41, 48, 49, 60, 67, 66, 70, 78, 87, 96, 101, 124, 128, 123, 136, 131, 143, 143, 138, 149, 146, 143, 147, 133, 138, 153, 148, 147, 145, 155, 158, 156, 156, 159, 159, 156, 157, 163, 158, 155, 163, 155, 148, 152, 149, 149, 139, 146, 138, 149, 149, 154, 156, 153, 158, 152, 156, 146, 145, 155, 165, 154, 140, 159, 151, 159, 159, 152, 157, 151, 154, 158, 139, 165, 159, 166, 165, 160, 134, 142, 146, 188, 177, 141, 152, 149, 151, 150, 161, 151, 148, 153, 156, 154, 156, 147, 156, 152, 158, 161, 135, 114, 117, 145, 168, 183, 203, 159, 148, 152, 152, 147, 150, 143, 155, 157, 146, 157, 148, 107, 106, 137, 163, 147, 149, 155, 147, 151, 156, 156, 156, 150, 150, 148, 149, 143, 146, 134, 158, 153, 146, 139, 150, 145, 152, 148, 149, 144, 141, 138, 166, 148, 149, 144, 144, 143, 153, 150, 139, 142, 139, 134, 143, 140, 140, 133, 140, 127, 133, 115, 146, 129, 130, 136, 106, 104, 125, 123, 132, 127, 125, 133, 132, 112, 122, 128, 123, 122, 137, 124, 113, 111, 106, 110, 109, 110, 111, 117, 114, 126, 116, 118, 123, 133, 128, 133, 141, 136, 135, 140, 131, 120, 113, 97, 88, 79, 72, 72, 76, 76, 85, 90, 94, 90, 114, 136, 147, 147, 168, 177, 171, 179, 190, 198, 206, 207, 211, 204, 211, 204, 204, 188, 181, 186, 177, 179, 154, 139, 110, 75, 60, 53, 52, 65, 48, 36, 38, 50, 54, 58, 60, 70, 71, 76, 87, 91, 109, 125, 132, 129, 142, 131, 138, 142, 142, 143, 146, 142, 151, 136, 146, 147, 143, 138, 151, 156, 158, 156, 159, 167, 153, 143, 160, 155, 152, 161, 154, 158, 156, 155, 149, 152, 138, 147, 141, 144, 154, 151, 155, 156, 159, 159, 150, 149, 142, 154, 159, 158, 150, 156, 158, 161, 157, 152, 166, 153, 156, 145, 146, 181, 163, 167, 170, 157, 105, 132, 156, 194, 215, 161, 139, 141, 149, 147, 162, 153, 157, 149, 144, 157, 156, 157, 157, 148, 156, 160, 137, 132, 116, 136, 156, 170, 175, 142, 142, 145, 149, 150, 152, 150, 153, 150, 151, 147, 149, 117, 86, 128, 137, 136, 146, 141, 138, 141, 156, 147, 133, 147, 182, 167, 148, 149, 140, 140, 148, 145, 140, 145, 147, 150, 154, 150, 153, 148, 142, 147, 135, 143, 149, 155, 143, 144, 150, 148, 140, 139, 138, 138, 139, 147, 142, 118, 136, 143, 135, 132, 124, 128, 127, 129, 122, 117, 123, 128, 128, 122, 127, 126, 123, 118, 119, 129, 128, 124, 127, 125, 119, 110, 104, 116, 111, 113, 118, 119, 112, 114, 118, 116, 117, 131, 136, 132, 133, 138, 131, 138, 132, 134, 117, 95, 93, 76, 72, 56, 67, 63, 63, 77, 90, 91, 100, 109, 132, 140, 158, 167, 176, 178, 187, 198, 196, 199, 200, 202, 205, 201, 195, 187, 192, 193, 174, 176, 175, 151, 102, 77, 58, 44, 46, 69, 59, 47, 41, 47, 59, 56, 64, 72, 63, 75, 76, 95, 95, 125, 125, 138, 136, 136, 140, 144, 144, 151, 148, 155, 149, 141, 148, 146, 137, 135, 143, 150, 158, 152, 146, 157, 162, 150, 155, 145, 158, 157, 151, 149, 146, 151, 148, 151, 150, 146, 138, 154, 158, 156, 160, 148, 160, 161, 159, 159, 125, 141, 157, 160, 159, 150, 158, 161, 157, 150, 146, 153, 163, 135, 156, 198, 181, 149, 174, 170, 96, 131, 148, 179, 221, 180, 132, 148, 156, 133, 153, 147, 145, 151, 149, 150, 157, 158, 153, 156, 149, 149, 143, 142, 130, 131, 139, 155, 145, 136, 141, 146, 149, 151, 151, 143, 148, 152, 147, 152, 151, 145, 137, 140, 138, 139, 141, 152, 143, 144, 142, 124, 98, 143, 181, 193, 148, 148, 140, 154, 163, 143, 150, 153, 143, 148, 150, 157, 151, 147, 145, 145, 135, 145, 148, 148, 148, 144, 147, 148, 137, 149, 143, 143, 139, 138, 146, 130, 142, 142, 130, 138, 119, 125, 125, 128, 130, 120, 116, 126, 131, 126, 121, 133, 131, 134, 131, 129, 121, 119, 127, 121, 126, 122, 117, 109, 113, 109, 108, 109, 108, 106, 106, 108, 119, 121, 113, 126, 122, 130, 122, 133, 131, 123, 118, 103, 92, 77, 64, 58, 62, 65, 60, 74, 78, 89, 94, 100, 132, 137, 152, 162, 172, 174, 176, 188, 198, 202, 192, 203, 201, 197, 203, 196, 187, 192, 180, 177, 175, 165, 123, 93, 70, 48, 50, 41, 45, 51, 49, 60, 68, 66, 54, 61, 58, 64, 68, 91, 94, 122, 135, 138, 135, 140, 140, 145, 144, 149, 142, 151, 153, 152, 141, 155, 151, 134, 142, 150, 155, 162, 145, 161, 160, 153, 155, 159, 151, 158, 154, 156, 150, 148, 150, 154, 141, 145, 147, 147, 155, 153, 148, 157, 155, 159, 158, 155, 144, 141, 155, 143, 155, 149, 158, 160, 157, 157, 147, 162, 156, 132, 160, 178, 179, 156, 154, 172, 78, 130, 144, 164, 204, 157, 130, 144, 141, 144, 143, 144, 148, 152, 143, 147, 149, 149, 147, 154, 157, 148, 155, 136, 152, 182, 137, 122, 139, 160, 172, 155, 151, 150, 150, 153, 148, 145, 146, 148, 153, 146, 136, 145, 142, 134, 144, 143, 142, 149, 145, 111, 91, 133, 171, 170, 136, 139, 149, 146, 155, 147, 146, 148, 148, 147, 135, 153, 149, 142, 138, 148, 146, 140, 144, 143, 140, 149, 150, 143, 132, 135, 142, 145, 140, 137, 139, 140, 143, 141, 135, 143, 138, 124, 131, 129, 130, 136, 127, 121, 127, 126, 132, 132, 132, 145, 141, 132, 125, 118, 118, 116, 118, 118, 108, 112, 107, 93, 104, 105, 94, 89, 95, 104, 106, 114, 126, 127, 129, 128, 133, 133, 132, 127, 117, 107, 81, 74, 68, 66, 68, 59, 55, 66, 76, 85, 90, 96, 109, 135, 143, 148, 166, 172, 179, 187, 189, 195, 197, 195, 195, 198, 197, 192, 196, 200, 193, 177, 169, 173, 145, 113, 89, 73, 63, 34, 45, 58, 53, 60, 66, 67, 54, 66, 59, 66, 73, 92, 97, 115, 135, 138, 142, 147, 144, 138, 142, 150, 157, 152, 155, 153, 147, 148, 154, 142, 149, 147, 161, 168, 139, 165, 159, 155, 154, 152, 167, 158, 147, 148, 150, 156, 160, 153, 138, 142, 147, 140, 152, 151, 141, 163, 156, 159, 158, 155, 157, 150, 156, 128, 133, 141, 158, 160, 150, 158, 151, 154, 162, 137, 160, 175, 163, 163, 167, 173, 94, 116, 143, 162, 163, 131, 144, 148, 145, 142, 138, 137, 148, 148, 143, 154, 148, 152, 148, 154, 152, 159, 148, 137, 145, 179, 134, 118, 130, 155, 198, 167, 147, 160, 148, 154, 150, 151, 146, 156, 132, 144, 152, 154, 147, 132, 142, 133, 143, 147, 146, 131, 102, 124, 160, 148, 133, 142, 145, 151, 150, 150, 140, 146, 147, 152, 150, 157, 151, 146, 140, 144, 147, 145, 147, 151, 136, 138, 144, 145, 145, 135, 139, 143, 141, 143, 146, 132, 140, 138, 127, 129, 138, 132, 127, 131, 127, 129, 131, 127, 136, 136, 133, 130, 139, 143, 134, 125, 116, 116, 110, 103, 118, 108, 108, 110, 102, 102, 94, 87, 66, 88, 91, 99, 111, 111, 118, 131, 141, 140, 141, 144, 143, 134, 113, 109, 94, 66, 68, 60, 66, 58, 49, 60, 71, 76, 84, 102, 102, 119, 133, 141, 151, 170, 172, 177, 186, 192, 194, 189, 192, 195, 191, 196, 189, 193, 203, 178, 177, 173, 152, 124, 117, 91, 69, 46, 53, 64, 65, 64, 68, 71, 67, 78, 64, 63, 69, 85, 99, 117, 139, 138, 143, 138, 135, 144, 145, 150, 155, 153, 156, 149, 144, 159, 160, 150, 159, 165, 165, 158, 152, 162, 161, 157, 157, 156, 165, 157, 156, 155, 155, 145, 157, 157, 153, 145, 150, 150, 152, 155, 157, 155, 151, 157, 156, 152, 152, 152, 152, 126, 131, 136, 149, 159, 148, 150, 171, 162, 148, 155, 165, 170, 159, 161, 170, 178, 133, 127, 129, 137, 125, 120, 142, 166, 147, 143, 140, 140, 133, 144, 136, 147, 157, 148, 150, 150, 150, 158, 157, 151, 149, 148, 109, 115, 128, 159, 184, 161, 139, 147, 142, 143, 147, 150, 147, 148, 133, 144, 137, 145, 152, 146, 143, 142, 141, 138, 141, 149, 142, 147, 140, 140, 133, 148, 155, 142, 141, 144, 148, 147, 126, 164, 159, 145, 154, 152, 143, 144, 143, 142, 143, 150, 144, 139, 144, 139, 138, 138, 141, 135, 142, 140, 137, 131, 146, 147, 138, 142, 138, 135, 134, 129, 123, 125, 122, 124, 121, 129, 145, 146, 142, 137, 135, 125, 119, 116, 113, 102, 114, 100, 105, 96, 83, 98, 106, 104, 93, 96, 94, 103, 118, 118, 123, 130, 141, 141, 148, 159, 149, 132, 126, 115, 103, 83, 74, 71, 60, 53, 58, 60, 59, 62, 82, 93, 101, 112, 133, 137, 134, 159, 165, 174, 181, 188, 185, 187, 189, 193, 195, 193, 196, 195, 204, 190, 181, 178, 166, 135, 126, 108, 87, 60, 53, 64, 62, 65, 70, 69, 73, 78, 58, 55, 61, 88, 97, 114, 127, 146, 140, 133, 130, 141, 148, 144, 153, 152, 157, 136, 150, 172, 166, 145, 179, 159, 158, 154, 158, 157, 159, 154, 148, 144, 157, 159, 158, 159, 161, 152, 163, 161, 163, 143, 152, 152, 147, 155, 155, 160, 160, 158, 149, 163, 158, 158, 136, 162, 145, 155, 154, 158, 135, 148, 174, 171, 154, 167, 162, 163, 165, 174, 176, 166, 147, 139, 123, 129, 136, 123, 138, 146, 126, 136, 122, 111, 124, 135, 138, 137, 147, 149, 156, 159, 159, 156, 156, 150, 148, 133, 117, 110, 126, 150, 172, 143, 148, 130, 145, 142, 131, 142, 142, 140, 145, 146, 144, 144, 140, 140, 147, 147, 145, 143, 140, 142, 144, 149, 151, 144, 135, 144, 143, 146, 143, 149, 144, 150, 133, 147, 148, 149, 147, 150, 145, 135, 161, 131, 140, 148, 160, 149, 136, 137, 138, 132, 140, 139, 134, 132, 138, 136, 128, 140, 139, 138, 137, 137, 139, 129, 121, 127, 132, 135, 125, 138, 151, 152, 146, 140, 139, 136, 121, 119, 111, 115, 100, 103, 101, 93, 82, 99, 100, 101, 85, 91, 91, 103, 125, 123, 121, 130, 140, 141, 149, 162, 148, 147, 135, 110, 102, 85, 75, 74, 69, 58, 59, 50, 65, 65, 75, 71, 96, 109, 126, 135, 133, 142, 158, 165, 171, 180, 179, 185, 186, 193, 188, 192, 193, 195, 203, 200, 190, 179, 166, 152, 118, 120, 96, 77, 72, 74, 52, 59, 65, 71, 77, 77, 55, 60, 62, 93, 101, 119, 136, 140, 140, 140, 142, 144, 145, 145, 146, 149, 155, 123, 143, 180, 172, 151, 159, 150, 167, 163, 153, 169, 164, 159, 146, 153, 164, 166, 154, 147, 158, 164, 155, 154, 153, 161, 148, 151, 149, 159, 157, 155, 169, 161, 158, 156, 160, 159, 157, 159, 158, 152, 150, 159, 141, 148, 164, 152, 145, 183, 163, 161, 165, 179, 174, 166, 151, 144, 104, 134, 142, 137, 142, 129, 127, 150, 112, 106, 86, 109, 127, 137, 133, 152, 147, 149, 153, 156, 146, 151, 143, 141, 132, 132, 118, 139, 143, 150, 141, 75, 144, 187, 130, 156, 151, 136, 143, 141, 144, 141, 135, 138, 142, 150, 147, 146, 145, 148, 138, 130, 146, 144, 141, 138, 145, 151, 155, 153, 147, 153, 145, 150, 143, 151, 153, 153, 143, 126, 145, 134, 138, 146, 150, 156, 142, 130, 136, 136, 139, 139, 125, 123, 136, 132, 128, 138, 140, 139, 136, 136, 139, 128, 127, 127, 134, 137, 129, 141, 154, 153, 144, 147, 152, 132, 130, 126, 128, 118, 106, 106, 106, 99, 97, 110, 104, 93, 65, 83, 92, 98, 117, 121, 130, 139, 136, 142, 142, 144, 163, 143, 139, 122, 107, 76, 77, 74, 51, 57, 62, 59, 53, 65, 73, 77, 78, 102, 126, 134, 139, 146, 137, 142, 157, 172, 171, 177, 181, 185, 187, 185, 192, 203, 204, 194, 196, 183, 176, 167, 126, 119, 103, 87, 81, 87, 60, 67, 67, 73, 83, 86, 71, 62, 72, 93, 97, 121, 135, 136, 139, 136, 145, 136, 129, 142, 150, 147, 150, 145, 150, 173, 154, 150, 168, 162, 159, 150, 158, 160, 172, 163, 160, 170, 164, 166, 161, 164, 159, 156, 152, 157, 157, 160, 152, 159, 155, 155, 153, 149, 157, 154, 160, 157, 163, 158, 170, 155, 164, 152, 148, 157, 156, 150, 156, 148, 161, 160, 180, 163, 158, 168, 166, 156, 144, 129, 131, 140, 144, 145, 133, 135, 118, 125, 80, 99, 111, 99, 126, 135, 136, 143, 142, 149, 150, 152, 149, 149, 145, 149, 139, 137, 135, 140, 143, 151, 136, 94, 115, 151, 124, 166, 178, 140, 141, 149, 134, 142, 135, 135, 128, 145, 140, 145, 142, 143, 140, 136, 137, 149, 170, 142, 135, 138, 141, 152, 147, 146, 132, 169, 151, 148, 146, 152, 149, 144, 140, 136, 135, 142, 143, 155, 135, 140, 142, 137, 146, 139, 131, 112, 110, 126, 138, 141, 135, 141, 138, 139, 129, 127, 130, 123, 131, 129, 135, 147, 143, 144, 160, 162, 154, 150, 142, 139, 138, 124, 119, 114, 114, 108, 109, 100, 103, 100, 92, 73, 84, 101, 113, 123, 131, 139, 144, 147, 151, 151, 164, 156, 146, 122, 105, 83, 65, 68, 57, 49, 57, 51, 51, 56, 61, 73, 70, 94, 115, 135, 134, 138, 133, 141, 137, 158, 173, 172, 169, 178, 184, 188, 196, 205, 203, 202, 196, 191, 180, 160, 140, 113, 105, 95, 93, 92, 79, 80, 68, 68, 77, 83, 69, 65, 74, 85, 95, 128, 140, 145, 140, 142, 149, 143, 136, 151, 150, 152, 149, 159, 157, 164, 155, 154, 167, 161, 167, 166, 157, 163, 166, 161, 167, 166, 173, 162, 158, 160, 161, 177, 152, 159, 160, 153, 156, 150, 148, 155, 147, 150, 156, 152, 157, 153, 157, 163, 167, 161, 164, 161, 165, 156, 165, 143, 151, 162, 148, 146, 193, 179, 159, 169, 179, 175, 151, 144, 138, 143, 134, 145, 138, 148, 135, 119, 113, 87, 99, 118, 134, 132, 152, 145, 138, 146, 146, 147, 152, 148, 135, 145, 151, 146, 142, 142, 115, 140, 146, 150, 129, 103, 123, 155, 176, 143, 145, 132, 126, 150, 166, 138, 137, 144, 138, 141, 145, 148, 129, 113, 133, 161, 203, 170, 131, 138, 140, 152, 146, 144, 147, 145, 144, 150, 144, 138, 153, 148, 144, 130, 130, 135, 121, 140, 137, 139, 142, 140, 138, 137, 138, 114, 101, 132, 139, 141, 119, 145, 120, 133, 149, 134, 133, 119, 128, 122, 140, 150, 155, 158, 162, 167, 160, 147, 143, 140, 144, 137, 132, 122, 124, 112, 120, 103, 99, 88, 83, 70, 86, 100, 117, 123, 129, 141, 147, 148, 160, 157, 156, 155, 144, 127, 111, 91, 80, 55, 44, 46, 57, 43, 52, 58, 56, 69, 69, 93, 108, 123, 129, 129, 133, 137, 136, 139, 142, 169, 173, 174, 185, 184, 192, 207, 202, 209, 201, 199, 187, 155, 148, 130, 114, 111, 96, 97, 95, 89, 74, 73, 72, 84, 75, 77, 77, 94, 106, 123, 140, 138, 144, 140, 147, 142, 139, 153, 148, 153, 155, 154, 156, 157, 158, 156, 165, 155, 169, 154, 151, 164, 166, 162, 162, 168, 173, 166, 163, 160, 159, 161, 155, 163, 158, 151, 152, 155, 155, 158, 147, 157, 157, 147, 159, 154, 152, 157, 159, 173, 167, 162, 165, 166, 158, 147, 155, 140, 136, 169, 188, 189, 165, 171, 174, 169, 157, 146, 147, 143, 148, 135, 148, 145, 136, 140, 117, 123, 119, 136, 134, 135, 145, 144, 149, 144, 145, 150, 143, 151, 161, 144, 146, 132, 136, 168, 147, 116, 143, 159, 144, 121, 129, 143, 151, 131, 136, 113, 119, 141, 172, 158, 137, 139, 143, 134, 136, 135, 102, 111, 117, 157, 197, 158, 128, 149, 139, 146, 158, 150, 149, 150, 148, 145, 150, 142, 149, 139, 144, 137, 134, 136, 128, 134, 136, 137, 141, 142, 141, 136, 137, 135, 129, 127, 136, 139, 106, 142, 134, 130, 125, 142, 132, 118, 127, 139, 138, 146, 140, 163, 166, 172, 164, 161, 158, 145, 135, 142, 138, 134, 128, 108, 119, 109, 107, 98, 77, 84, 92, 93, 97, 113, 126, 141, 152, 158, 166, 157, 154, 156, 146, 120, 103, 83, 78, 55, 52, 47, 61, 49, 57, 66, 45, 50, 66, 81, 109, 109, 112, 126, 124, 129, 141, 137, 144, 140, 160, 165, 168, 175, 183, 195, 202, 203, 205, 195, 182, 164, 147, 141, 105, 97, 104, 97, 91, 91, 75, 67, 73, 76, 78, 78, 84, 98, 101, 140, 130, 155, 137, 150, 144, 140, 140, 143, 153, 149, 150, 155, 159, 161, 159, 157, 165, 156, 168, 165, 163, 157, 167, 169, 159, 166, 173, 156, 165, 163, 162, 157, 156, 153, 150, 149, 159, 158, 153, 159, 149, 153, 160, 145, 155, 168, 155, 156, 168, 158, 188, 160, 156, 169, 161, 153, 150, 142, 122, 164, 173, 188, 170, 165, 167, 158, 150, 150, 146, 148, 150, 130, 151, 146, 138, 138, 144, 133, 142, 133, 136, 150, 137, 138, 144, 139, 150, 134, 123, 144, 182, 155, 127, 103, 130, 170, 172, 132, 133, 143, 141, 138, 138, 133, 135, 131, 129, 106, 118, 125, 177, 169, 120, 129, 139, 140, 140, 130, 95, 94, 97, 150, 174, 134, 115, 127, 137, 139, 152, 151, 149, 142, 150, 149, 147, 149, 140, 145, 137, 130, 134, 127, 126, 124, 130, 134, 131, 135, 135, 133, 130, 131, 125, 124, 136, 133, 127, 119, 116, 123, 124, 132, 138, 118, 121, 140, 134, 150, 149, 159, 164, 164, 163, 159, 164, 152, 143, 145, 145, 143, 147, 119, 118, 123, 112, 101, 86, 79, 85, 85, 99, 110, 116, 133, 145, 164, 164, 159, 151, 148, 142, 119, 108, 99, 84, 73, 75, 56, 57, 54, 61, 63, 50, 45, 65, 79, 100, 124, 117, 125, 114, 134, 131, 133, 137, 132, 129, 151, 149, 167, 166, 173, 204, 203, 203, 188, 178, 164, 152, 140, 117, 110, 106, 100, 94, 94, 82, 74, 71, 78, 81, 86, 88, 100, 108, 139, 136, 145, 143, 149, 141, 149, 148, 142, 151, 150, 153, 153, 146, 157, 157, 166, 160, 162, 166, 165, 158, 161, 161, 159, 158, 165, 167, 164, 166, 165, 159, 161, 171, 160, 154, 152, 161, 162, 156, 156, 154, 152, 166, 143, 146, 167, 165, 162, 173, 106, 199, 185, 157, 162, 165, 157, 158, 148, 130, 152, 166, 168, 161, 173, 177, 160, 138, 155, 156, 151, 148, 143, 148, 147, 149, 146, 144, 149, 137, 135, 141, 124, 170, 133, 147, 142, 139, 129, 115, 143, 156, 143, 123, 99, 114, 146, 178, 134, 133, 136, 129, 134, 132, 130, 132, 127, 124, 97, 105, 139, 167, 154, 123, 127, 136, 138, 142, 128, 98, 112, 103, 144, 138, 114, 150, 151, 133, 154, 145, 144, 147, 141, 140, 143, 143, 140, 143, 141, 143, 127, 139, 132, 129, 128, 132, 130, 129, 140, 136, 133, 126, 122, 123, 120, 116, 107, 114, 122, 117, 126, 122, 118, 128, 136, 126, 142, 136, 144, 157, 156, 159, 159, 157, 156, 160, 157, 141, 137, 144, 151, 144, 129, 123, 120, 100, 105, 99, 73, 73, 78, 92, 102, 105, 123, 146, 157, 167, 167, 158, 144, 143, 124, 109, 112, 97, 83, 78, 80, 62, 59, 74, 57, 54, 55, 66, 86, 105, 126, 120, 117, 120, 129, 129, 124, 126, 138, 131, 134, 140, 159, 166, 168, 193, 197, 194, 192, 180, 168, 152, 142, 139, 120, 108, 105, 101, 102, 90, 91, 84, 80, 89, 87, 102, 102, 116, 132, 147, 138, 147, 144, 153, 150, 149, 150, 149, 150, 155, 154, 156, 158, 154, 165, 170, 161, 155, 168, 153, 174, 162, 160, 159, 165, 172, 165, 166, 175, 166, 155, 165, 160, 159, 157, 161, 160, 153, 158, 155, 151, 159, 156, 149, 161, 155, 159, 171, 126, 176, 171, 157, 161, 159, 158, 167, 170, 149, 144, 164, 161, 163, 161, 170, 161, 151, 156, 153, 154, 148, 148, 140, 152, 157, 141, 153, 147, 149, 138, 145, 106, 165, 144, 144, 147, 142, 137, 111, 131, 135, 127, 131, 100, 119, 135, 148, 144, 134, 136, 137, 108, 131, 144, 128, 131, 120, 95, 90, 134, 194, 164, 129, 121, 133, 128, 121, 151, 135, 123, 126, 133, 122, 121, 138, 160, 147, 150, 151, 144, 138, 150, 161, 145, 146, 144, 138, 134, 140, 135, 138, 129, 129, 130, 123, 123, 119, 128, 132, 126, 140, 132, 123, 104, 87, 76, 93, 135, 146, 146, 129, 112, 129, 133, 132, 138, 141, 153, 146, 153, 156, 161, 161, 163, 167, 157, 154, 142, 122, 143, 145, 136, 121, 127, 107, 93, 98, 73, 63, 69, 87, 94, 106, 112, 141, 147, 164, 166, 155, 144, 142, 129, 113, 104, 98, 94, 84, 81, 68, 62, 65, 66, 61, 57, 67, 76, 99, 115, 111, 123, 127, 131, 131, 118, 123, 137, 132, 130, 129, 144, 163, 169, 189, 187, 191, 183, 182, 171, 159, 144, 147, 121, 114, 110, 103, 114, 112, 108, 89, 85, 83, 86, 95, 109, 115, 140, 134, 133, 153, 148, 151, 150, 148, 150, 147, 151, 152, 155, 158, 160, 164, 167, 165, 167, 164, 163, 150, 173, 168, 163, 171, 168, 169, 170, 171, 179, 164, 164, 165, 158, 158, 156, 161, 155, 146, 166, 158, 158, 155, 158, 157, 159, 150, 150, 158, 166, 167, 166, 157, 166, 152, 149, 161, 156, 156, 164, 160, 164, 141, 173, 168, 167, 140, 153, 141, 159, 149, 148, 147, 118, 156, 156, 146, 140, 135, 148, 144, 143, 138, 133, 144, 140, 150, 132, 133, 153, 134, 136, 133, 130, 129, 133, 123, 133, 125, 131, 132, 94, 127, 165, 160, 130, 119, 82, 82, 125, 194, 205, 163, 130, 131, 126, 135, 129, 138, 137, 140, 141, 137, 126, 138, 149, 139, 148, 149, 138, 130, 149, 165, 150, 144, 133, 137, 131, 133, 139, 138, 119, 124, 161, 126, 120, 120, 133, 127, 125, 132, 135, 136, 99, 60, 58, 96, 148, 172, 184, 156, 124, 127, 126, 117, 134, 134, 150, 151, 153, 152, 157, 166, 161, 168, 159, 155, 150, 143, 147, 143, 152, 133, 110, 119, 119, 93, 72, 81, 68, 79, 85, 100, 112, 134, 149, 160, 164, 157, 138, 122, 124, 111, 113, 110, 102, 91, 86, 82, 66, 65, 54, 57, 61, 67, 72, 83, 117, 125, 132, 123, 124, 133, 123, 134, 133, 127, 132, 129, 137, 160, 163, 177, 189, 187, 183, 170, 167, 159, 147, 133, 94, 103, 96, 111, 109, 104, 103, 101, 92, 90, 87, 101, 101, 116, 135, 135, 140, 143, 148, 150, 149, 149, 152, 149, 159, 152, 150, 153, 156, 159, 160, 164, 166, 172, 157, 161, 165, 171, 165, 170, 167, 166, 173, 171, 172, 134, 170, 199, 153, 164, 167, 165, 153, 151, 158, 158, 160, 162, 160, 153, 154, 155, 152, 156, 162, 166, 163, 162, 161, 157, 152, 165, 142, 148, 170, 154, 160, 147, 175, 165, 176, 152, 150, 146, 141, 154, 147, 158, 133, 140, 143, 143, 149, 140, 151, 140, 151, 141, 141, 148, 138, 150, 144, 145, 146, 144, 145, 146, 123, 121, 156, 153, 150, 136, 136, 134, 87, 93, 143, 162, 130, 110, 84, 89, 128, 179, 210, 204, 148, 127, 130, 138, 138, 143, 142, 140, 143, 142, 136, 139, 141, 137, 144, 145, 144, 137, 149, 148, 132, 136, 147, 128, 138, 142, 144, 135, 117, 108, 154, 133, 125, 124, 126, 124, 124, 124, 134, 119, 74, 48, 41, 97, 157, 184, 203, 194, 135, 129, 118, 129, 137, 145, 145, 154, 156, 154, 145, 163, 165, 163, 162, 153, 148, 138, 151, 150, 145, 131, 121, 120, 112, 102, 72, 68, 76, 78, 75, 105, 115, 129, 144, 144, 155, 156, 140, 125, 117, 108, 111, 112, 115, 108, 103, 92, 73, 73, 62, 64, 59, 65, 77, 91, 117, 135, 127, 123, 116, 125, 122, 128, 132, 135, 136, 133, 136, 138, 159, 172, 176, 183, 178, 177, 171, 159, 156, 135, 123, 116, 113, 118, 121, 118, 106, 103, 92, 99, 105, 107, 89, 121, 134, 140, 141, 154, 143, 152, 151, 147, 131, 145, 171, 151, 153, 158, 155, 155, 151, 160, 185, 200, 168, 163, 167, 169, 172, 159, 168, 169, 172, 170, 165, 126, 159, 199, 167, 146, 168, 204, 162, 165, 157, 160, 159, 158, 152, 154, 158, 161, 164, 157, 143, 166, 143, 170, 165, 160, 160, 158, 157, 156, 163, 166, 156, 172, 161, 161, 172, 151, 148, 150, 139, 148, 149, 149, 154, 153, 135, 135, 150, 149, 153, 151, 151, 148, 150, 143, 145, 160, 149, 145, 146, 144, 145, 140, 116, 112, 131, 154, 150, 140, 132, 139, 115, 97, 134, 130, 110, 98, 80, 88, 122, 153, 182, 203, 161, 130, 137, 141, 138, 145, 147, 142, 143, 148, 151, 144, 144, 144, 154, 150, 138, 140, 148, 139, 132, 132, 151, 138, 139, 136, 141, 132, 127, 124, 124, 123, 129, 123, 123, 137, 119, 121, 141, 103, 65, 40, 19, 74, 153, 188, 208, 214, 149, 120, 123, 127, 133, 144, 156, 150, 154, 145, 153, 150, 160, 172, 174, 154, 141, 143, 144, 146, 145, 133, 132, 121, 112, 99, 87, 82, 82, 82, 78, 97, 105, 120, 142, 150, 150, 145, 128, 119, 106, 112, 109, 108, 118, 109, 102, 90, 75, 68, 61, 57, 64, 66, 75, 88, 114, 131, 132, 131, 123, 124, 124, 126, 127, 132, 141, 139, 134, 131, 141, 165, 163, 183, 179, 170, 167, 166, 145, 147, 141, 137, 121, 121, 125, 124, 118, 98, 92, 100, 112, 114, 108, 134, 143, 140, 137, 166, 146, 149, 157, 152, 139, 144, 156, 148, 151, 158, 160, 160, 119, 145, 181, 205, 188, 165, 159, 162, 162, 165, 163, 170, 174, 161, 161, 163, 165, 168, 168, 130, 161, 201, 173, 165, 160, 158, 155, 160, 157, 155, 156, 157, 166, 161, 158, 165, 155, 163, 160, 156, 155, 146, 155, 155, 163, 165, 157, 180, 163, 166, 163, 143, 141, 145, 144, 145, 147, 147, 132, 141, 163, 154, 140, 145, 154, 153, 146, 150, 145, 138, 136, 141, 153, 150, 143, 150, 143, 142, 133, 122, 137, 145, 144, 133, 132, 131, 147, 122, 135, 127, 114, 76, 83, 86, 106, 156, 172, 189, 148, 126, 131, 136, 139, 141, 136, 139, 139, 147, 146, 135, 118, 144, 162, 151, 147, 142, 143, 141, 147, 135, 137, 154, 143, 137, 134, 134, 135, 140, 134, 132, 125, 128, 115, 141, 122, 118, 146, 118, 63, 25, 22, 80, 136, 168, 195, 198, 142, 124, 128, 136, 137, 137, 146, 146, 151, 150, 160, 162, 171, 173, 173, 153, 131, 144, 148, 148, 148, 127, 130, 119, 115, 98, 83, 84, 73, 77, 81, 89, 107, 115, 132, 138, 140, 139, 133, 124, 113, 115, 111, 118, 111, 96, 99, 80, 77, 78, 60, 53, 74, 75, 78, 85, 118, 127, 128, 121, 123, 125, 126, 123, 124, 126, 143, 136, 137, 129, 135, 150, 150, 176, 171, 164, 159, 156, 150, 154, 143, 142, 122, 124, 122, 127, 121, 101, 93, 104, 124, 123, 128, 137, 142, 139, 141, 149, 139, 148, 156, 153, 146, 158, 145, 156, 170, 161, 139, 170, 149, 137, 165, 197, 183, 163, 173, 177, 162, 165, 169, 167, 163, 163, 163, 165, 172, 163, 172, 158, 141, 172, 164, 166, 158, 157, 147, 156, 157, 165, 151, 150, 155, 159, 167, 159, 158, 163, 157, 160, 155, 162, 149, 158, 160, 160, 142, 186, 169, 173, 164, 134, 152, 148, 138, 149, 149, 153, 143, 109, 154, 164, 146, 152, 148, 143, 139, 149, 141, 142, 147, 142, 144, 144, 144, 152, 143, 143, 138, 122, 127, 125, 135, 142, 134, 148, 133, 143, 155, 136, 126, 104, 83, 66, 86, 124, 145, 162, 139, 129, 130, 142, 142, 143, 138, 140, 147, 149, 148, 138, 122, 147, 150, 141, 139, 167, 139, 127, 152, 137, 122, 153, 148, 126, 128, 133, 129, 134, 132, 134, 130, 132, 124, 130, 124, 127, 139, 128, 85, 47, 56, 95, 129, 155, 175, 163, 116, 125, 123, 125, 125, 144, 143, 145, 141, 134, 154, 162, 172, 177, 168, 158, 131, 137, 145, 148, 157, 140, 123, 120, 118, 93, 75, 89, 90, 83, 79, 91, 110, 129, 118, 137, 142, 133, 139, 126, 116, 108, 123, 121, 114, 106, 95, 86, 79, 74, 65, 70, 72, 79, 81, 95, 115, 121, 126, 127, 124, 126, 120, 125, 128, 124, 143, 130, 135, 121, 129, 145, 153, 166, 163, 155, 148, 148, 148, 156, 151, 146, 129, 124, 115, 124, 121, 107, 105, 115, 129, 123, 132, 139, 143, 149, 146, 149, 144, 144, 153, 158, 152, 155, 144, 150, 175, 165, 149, 161, 149, 138, 163, 176, 166, 158, 171, 167, 171, 159, 158, 168, 158, 160, 165, 169, 167, 167, 169, 167, 173, 165, 151, 169, 179, 159, 155, 151, 141, 175, 185, 148, 157, 153, 161, 160, 136, 149, 163, 161, 159, 160, 156, 151, 147, 164, 164, 165, 162, 173, 155, 145, 147, 151, 154, 155, 152, 146, 145, 124, 137, 149, 142, 157, 143, 132, 127, 148, 140, 149, 138, 139, 145, 143, 140, 145, 150, 146, 136, 145, 139, 142, 136, 143, 138, 132, 136, 147, 161, 139, 145, 145, 126, 102, 94, 108, 128, 138, 136, 135, 131, 133, 144, 143, 137, 130, 136, 149, 141, 133, 141, 145, 121, 109, 145, 165, 137, 124, 157, 150, 130, 133, 130, 120, 128, 131, 132, 133, 138, 132, 133, 132, 128, 124, 129, 129, 126, 130, 104, 70, 60, 82, 103, 127, 135, 111, 104, 121, 131, 125, 122, 138, 136, 133, 132, 136, 146, 157, 163, 174, 166, 148, 135, 135, 132, 132, 152, 139, 112, 123, 114, 103, 96, 91, 94, 84, 75, 96, 107, 119, 115, 131, 149, 142, 127, 124, 91, 95, 111, 124, 115, 97, 94, 90, 87, 77, 77, 77, 77, 76, 90, 96, 113, 115, 121, 122, 128, 124, 122, 130, 126, 129, 133, 128, 130, 131, 141, 147, 152, 146, 154, 150, 142, 140, 146, 146, 150, 145, 143, 137, 128, 124, 117, 121, 116, 120, 136, 136, 150, 145, 146, 152, 147, 150, 151, 150, 119, 163, 191, 153, 160, 159, 162, 165, 161, 165, 159, 162, 154, 156, 158, 162, 160, 166, 171, 163, 164, 157, 168, 163, 159, 167, 168, 158, 171, 164, 165, 165, 165, 159, 200, 158, 160, 146, 132, 166, 186, 155, 158, 156, 153, 158, 130, 152, 157, 156, 158, 157, 151, 149, 133, 153, 157, 158, 161, 168, 172, 141, 150, 146, 142, 151, 150, 145, 150, 145, 146, 153, 136, 146, 150, 143, 134, 150, 141, 143, 146, 139, 137, 141, 144, 139, 147, 127, 141, 141, 149, 144, 142, 139, 133, 127, 137, 124, 149, 138, 144, 139, 129, 133, 126, 108, 127, 125, 135, 136, 135, 138, 135, 137, 133, 134, 139, 146, 137, 139, 139, 143, 144, 107, 160, 153, 126, 120, 152, 164, 149, 125, 128, 123, 128, 130, 131, 127, 127, 130, 126, 123, 118, 115, 122, 119, 126, 126, 119, 105, 93, 94, 96, 103, 105, 95, 95, 128, 130, 126, 129, 133, 133, 130, 130, 135, 149, 154, 153, 152, 165, 149, 135, 134, 124, 124, 133, 117, 87, 120, 120, 115, 110, 96, 96, 84, 84, 89, 109, 130, 93, 122, 143, 126, 127, 122, 115, 106, 113, 118, 112, 103, 101, 86, 76, 71, 77, 78, 86, 79, 88, 99, 111, 115, 122, 130, 128, 125, 126, 127, 126, 130, 131, 134, 134, 127, 140, 147, 147, 138, 136, 138, 141, 134, 146, 151, 143, 142, 147, 137, 129, 130, 130, 125, 125, 129, 145, 143, 147, 149, 144, 148, 149, 152, 155, 155, 101, 146, 191, 147, 150, 163, 154, 158, 160, 162, 158, 159, 161, 156, 165, 173, 159, 164, 171, 156, 173, 160, 159, 162, 169, 156, 164, 171, 169, 162, 163, 166, 158, 155, 166, 160, 165, 164, 131, 155, 156, 156, 164, 165, 151, 163, 156, 160, 163, 153, 154, 154, 159, 150, 150, 159, 159, 160, 151, 155, 156, 140, 159, 151, 146, 145, 146, 150, 150, 144, 138, 141, 135, 145, 143, 143, 143, 140, 135, 132, 138, 142, 138, 131, 139, 134, 145, 121, 136, 145, 143, 142, 140, 142, 135, 132, 113, 136, 148, 140, 144, 134, 131, 133, 138, 127, 132, 130, 137, 136, 129, 138, 134, 128, 131, 135, 130, 139, 140, 146, 136, 149, 143, 112, 141, 137, 106, 119, 161, 171, 164, 121, 113, 111, 120, 122, 128, 131, 127, 125, 126, 129, 117, 119, 104, 109, 119, 115, 125, 128, 114, 93, 108, 91, 89, 121, 116, 126, 136, 129, 128, 129, 132, 124, 128, 126, 146, 144, 149, 152, 160, 152, 141, 132, 124, 122, 108, 108, 114, 123, 118, 117, 114, 104, 96, 103, 87, 91, 103, 120, 104, 105, 126, 130, 121, 107, 107, 117, 113, 122, 117, 99, 94, 89, 74, 77, 86, 85, 84, 94, 93, 105, 115, 117, 127, 132, 122, 119, 133, 122, 121, 130, 137, 132, 133, 136, 138, 148, 144, 138, 128, 132, 138, 135, 142, 158, 142, 146, 145, 137, 136, 116, 132, 132, 132, 135, 147, 145, 141, 152, 147, 140, 146, 158, 148, 160, 132, 136, 169, 145, 155, 155, 156, 160, 149, 154, 162, 159, 161, 169, 165, 168, 162, 156, 164, 166, 158, 161, 165, 172, 164, 162, 160, 171, 167, 162, 162, 167, 163, 159, 169, 153, 152, 180, 166, 154, 162, 156, 166, 169, 164, 153, 160, 160, 162, 149, 149, 151, 161, 161, 150, 155, 164, 153, 162, 150, 158, 147, 146, 148, 149, 145, 159, 142, 148, 150, 150, 144, 124, 155, 139, 144, 142, 146, 149, 133, 142, 152, 144, 142, 147, 155, 152, 152, 136, 146, 144, 132, 132, 153, 149, 135, 111, 135, 135, 135, 143, 137, 129, 124, 137, 140, 116, 133, 144, 137, 135, 127, 118, 128, 123, 140, 142, 134, 136, 136, 127, 145, 138, 117, 138, 120, 92, 118, 167, 167, 157, 128, 108, 107, 106, 110, 122, 120, 122, 111, 119, 126, 116, 114, 111, 103, 104, 106, 116, 116, 114, 92, 104, 111, 128, 128, 121, 124, 136, 125, 140, 137, 124, 117, 124, 125, 140, 145, 147, 150, 159, 149, 144, 138, 134, 120, 104, 105, 127, 125, 110, 107, 111, 104, 105, 100, 97, 105, 107, 102, 92, 109, 125, 136, 128, 118, 99, 89, 111, 122, 122, 104, 96, 89, 84, 87, 83, 87, 92, 102, 101, 117, 118, 114, 123, 125, 122, 124, 120, 117, 118, 126, 136, 135, 132, 132, 126, 143, 144, 136, 123, 122, 131, 128, 130, 137, 146, 149, 153, 142, 135, 128, 132, 139, 145, 144, 149, 148, 148, 142, 152, 142, 148, 153, 149, 159, 148, 149, 151, 149, 154, 150, 160, 159, 150, 151, 165, 159, 160, 171, 152, 161, 161, 161, 172, 160, 169, 162, 156, 173, 158, 163, 162, 167, 164, 165, 167, 165, 169, 159, 163, 150, 146, 166, 165, 135, 190, 169, 152, 165, 160, 161, 161, 161, 161, 158, 152, 157, 157, 156, 147, 159, 150, 151, 154, 157, 165, 141, 155, 152, 152, 153, 150, 141, 146, 155, 140, 140, 143, 142, 143, 145, 145, 141, 154, 143, 144, 149, 147, 138, 137, 142, 163, 150, 143, 144, 138, 143, 128, 150, 139, 142, 137, 126, 132, 136, 138, 131, 134, 120, 133, 132, 124, 128, 132, 127, 130, 125, 128, 121, 137, 135, 134, 128, 141, 125, 123, 144, 130, 117, 156, 115, 99, 112, 157, 166, 167, 164, 150, 135, 122, 124, 119, 127, 121, 117, 116, 116, 115, 106, 105, 99, 99, 108, 108, 114, 101, 107, 103, 112, 118, 125, 130, 133, 130, 129, 129, 136, 123, 122, 113, 104, 106, 139, 140, 143, 152, 152, 139, 120, 129, 123, 109, 104, 119, 121, 116, 108, 98, 104, 97, 97, 102, 110, 112, 114, 89, 97, 119, 126, 127, 124, 98, 87, 113, 121, 129, 116, 96, 95, 89, 93, 86, 94, 98, 109, 122, 122, 120, 123, 120, 127, 124, 126, 119, 120, 128, 129, 129, 127, 131, 132, 138, 144, 145, 133, 124, 120, 129, 119, 126, 128, 143, 142, 150, 144, 138, 125, 125, 138, 145, 140, 149, 151, 147, 150, 149, 148, 148, 154, 155, 153, 159, 161, 152, 154, 144, 151, 152, 156, 157, 153, 153, 152, 163, 165, 149, 165, 156, 141, 184, 159, 161, 161, 161, 167, 161, 165, 158, 166, 161, 162, 165, 159, 180, 165, 157, 155, 145, 174, 145, 112, 195, 192, 159, 150, 159, 158, 158, 155, 156, 153, 161, 138, 162, 153, 148, 151, 151, 150, 155, 162, 167, 150, 153, 137, 154, 146, 140, 143, 153, 143, 146, 142, 135, 148, 143, 142, 141, 136, 152, 149, 146, 152, 139, 128, 135, 127, 150, 156, 141, 141, 142, 140, 146, 135, 127, 146, 158, 137, 137, 142, 133, 131, 141, 139, 131, 126, 132, 125, 135, 128, 132, 120, 120, 108, 136, 115, 106, 142, 187, 164, 128, 137, 118, 141, 151, 114, 101, 92, 147, 161, 165, 185, 181, 155, 118, 101, 118, 126, 124, 111, 114, 117, 112, 104, 104, 106, 96, 100, 104, 103, 107, 107, 124, 156, 118, 125, 134, 124, 130, 138, 125, 128, 129, 120, 111, 92, 63, 111, 150, 151, 140, 140, 138, 132, 129, 123, 116, 108, 100, 117, 113, 96, 103, 109, 109, 95, 103, 118, 112, 94, 82, 91, 106, 115, 126, 126, 120, 113, 117, 118, 118, 106, 108, 102, 95, 98, 94, 100, 114, 117, 132, 130, 116, 118, 119, 124, 126, 134, 117, 121, 128, 119, 122, 124, 134, 123, 126, 148, 163, 131, 113, 105, 113, 109, 119, 117, 129, 142, 142, 141, 141, 117, 139, 137, 142, 150, 147, 154, 143, 154, 150, 146, 147, 156, 147, 155, 158, 154, 148, 157, 154, 146, 161, 151, 163, 163, 155, 158, 143, 160, 158, 162, 154, 153, 161, 161, 162, 166, 156, 152, 203, 167, 164, 153, 179, 161, 166, 166, 171, 162, 157, 164, 158, 159, 161, 133, 170, 161, 172, 160, 165, 154, 160, 157, 157, 152, 166, 157, 155, 148, 161, 156, 147, 157, 144, 166, 162, 148, 146, 141, 153, 151, 148, 150, 152, 139, 131, 149, 142, 140, 140, 134, 147, 131, 141, 140, 148, 146, 144, 134, 144, 131, 142, 156, 138, 134, 146, 141, 141, 149, 137, 128, 139, 127, 135, 142, 137, 123, 129, 140, 131, 128, 126, 125, 128, 122, 107, 123, 186, 146, 116, 83, 86, 138, 192, 202, 127, 123, 127, 131, 138, 105, 97, 91, 106, 124, 147, 164, 179, 176, 138, 104, 101, 113, 121, 114, 110, 110, 113, 111, 114, 115, 110, 107, 120, 118, 115, 100, 95, 139, 141, 129, 124, 112, 116, 133, 127, 126, 124, 125, 126, 100, 82, 125, 156, 156, 139, 133, 129, 123, 116, 122, 114, 116, 99, 109, 107, 94, 91, 99, 102, 111, 118, 131, 118, 100, 79, 85, 100, 121, 128, 138, 129, 122, 128, 124, 112, 109, 107, 103, 98, 94, 103, 113, 120, 131, 141, 137, 125, 118, 123, 120, 123, 130, 122, 119, 123, 124, 126, 124, 126, 109, 111, 152, 178, 145, 120, 99, 98, 97, 112, 113, 119, 129, 144, 137, 143, 140, 141, 141, 144, 149, 148, 145, 151, 157, 151, 147, 151, 155, 150, 157, 152, 151, 152, 154, 158, 150, 149, 145, 160, 152, 158, 178, 149, 151, 156, 153, 153, 160, 166, 158, 163, 166, 157, 136, 195, 169, 163, 152, 172, 165, 164, 167, 171, 167, 158, 165, 162, 158, 164, 161, 156, 155, 163, 157, 167, 154, 165, 160, 152, 162, 155, 152, 155, 158, 162, 153, 146, 157, 152, 165, 157, 142, 142, 146, 147, 144, 146, 142, 141, 142, 144, 146, 145, 136, 133, 144, 139, 157, 138, 141, 144, 136, 145, 131, 148, 144, 121, 147, 144, 140, 147, 142, 141, 140, 145, 138, 134, 136, 128, 135, 130, 130, 132, 132, 129, 127, 123, 121, 129, 109, 72, 85, 184, 175, 119, 73, 74, 136, 173, 197, 135, 132, 131, 127, 142, 122, 117, 100, 90, 118, 127, 119, 170, 199, 183, 158, 115, 93, 107, 120, 114, 114, 107, 116, 115, 111, 113, 116, 121, 124, 120, 117, 101, 122, 138, 126, 123, 120, 107, 117, 113, 129, 128, 130, 123, 98, 84, 107, 132, 143, 138, 129, 126, 123, 110, 116, 113, 112, 116, 106, 119, 112, 109, 103, 100, 117, 122, 126, 122, 103, 99, 90, 85, 100, 123, 137, 136, 129, 123, 120, 114, 109, 102, 110, 105, 102, 104, 107, 118, 129, 149, 139, 123, 116, 118, 121, 117, 119, 123, 120, 119, 133, 126, 116, 121, 121, 109, 146, 157, 143, 129, 118, 110, 98, 98, 96, 120, 123, 135, 137, 146, 146, 134, 145, 144, 153, 146, 140, 141, 149, 153, 140, 158, 150, 147, 157, 152, 154, 153, 152, 151, 154, 150, 144, 151, 128, 159, 183, 172, 155, 151, 155, 159, 166, 165, 164, 161, 165, 166, 158, 164, 160, 161, 156, 167, 172, 161, 166, 172, 164, 163, 158, 160, 166, 154, 166, 156, 157, 159, 159, 163, 158, 156, 156, 161, 160, 158, 155, 152, 155, 149, 142, 152, 151, 167, 156, 156, 155, 147, 142, 145, 150, 143, 139, 149, 143, 143, 151, 138, 140, 139, 143, 138, 147, 140, 153, 150, 132, 135, 142, 131, 136, 125, 140, 146, 143, 141, 129, 132, 142, 136, 129, 142, 139, 143, 128, 128, 125, 130, 126, 120, 128, 104, 132, 145, 123, 104, 77, 148, 138, 131, 99, 79, 129, 156, 158, 124, 131, 138, 136, 135, 124, 124, 136, 94, 122, 94, 67, 124, 187, 198, 208, 178, 113, 108, 108, 111, 112, 105, 116, 126, 121, 111, 116, 119, 122, 126, 131, 117, 124, 128, 123, 128, 133, 121, 125, 116, 130, 121, 128, 123, 106, 91, 107, 121, 116, 119, 123, 116, 128, 112, 110, 93, 102, 107, 103, 111, 118, 117, 115, 101, 108, 119, 136, 133, 97, 109, 91, 91, 85, 108, 127, 139, 133, 128, 118, 106, 105, 100, 106, 121, 114, 111, 107, 126, 133, 145, 137, 129, 119, 118, 122, 125, 131, 132, 121, 123, 125, 128, 123, 126, 127, 131, 139, 152, 140, 137, 125, 111, 118, 109, 107, 117, 123, 133, 137, 139, 140, 145, 148, 148, 139, 146, 152, 150, 148, 153, 147, 147, 159, 159, 155, 157, 157, 156, 155, 150, 153, 153, 151, 147, 133, 150, 168, 171, 164, 150, 165, 157, 164, 169, 159, 165, 155, 167, 171, 167, 163, 154, 158, 165, 165, 168, 171, 164, 167, 160, 159, 157, 156, 161, 163, 156, 165, 159, 157, 160, 151, 156, 157, 160, 160, 161, 158, 155, 150, 140, 155, 156, 148, 154, 155, 153, 143, 142, 142, 135, 144, 140, 148, 147, 136, 149, 141, 122, 163, 147, 138, 149, 142, 130, 150, 144, 143, 138, 145, 138, 130, 129, 125, 124, 143, 152, 112, 118, 120, 122, 143, 135, 134, 143, 127, 126, 129, 135, 123, 131, 117, 97, 151, 175, 131, 138, 123, 133, 128, 136, 125, 96, 111, 138, 124, 125, 131, 134, 140, 132, 124, 130, 144, 105, 110, 80, 62, 89, 131, 168, 199, 203, 158, 115, 101, 122, 123, 123, 110, 124, 123, 129, 121, 125, 126, 125, 122, 123, 114, 149, 130, 125, 133, 124, 117, 115, 126, 121, 118, 120, 119, 109, 113, 107, 117, 114, 106, 110, 119, 112, 108, 107, 94, 98, 103, 112, 121, 116, 114, 123, 119, 122, 139, 135, 116, 100, 101, 92, 91, 98, 117, 132, 133, 130, 117, 107, 91, 108, 105, 119, 116, 124, 116, 122, 135, 141, 139, 127, 122, 130, 123, 135, 129, 125, 131, 134, 124, 122, 122, 128, 133, 136, 155, 155, 137, 139, 135, 124, 125, 124, 116, 113, 119, 125, 134, 142, 145, 155, 144, 147, 150, 145, 144, 153, 147, 150, 157, 141, 159, 154, 154, 156, 155, 153, 154, 155, 155, 152, 158, 154, 153, 151, 161, 152, 156, 155, 163, 161, 160, 166, 161, 158, 154, 165, 161, 175, 167, 151, 172, 167, 165, 161, 169, 166, 163, 162, 165, 157, 159, 166, 169, 158, 173, 164, 160, 168, 158, 151, 162, 157, 159, 163, 158, 149, 158, 151, 158, 151, 152, 151, 151, 161, 144, 131, 154, 143, 142, 143, 143, 144, 129, 138, 146, 126, 149, 153, 139, 148, 139, 143, 146, 134, 132, 138, 135, 138, 138, 134, 149, 122, 125, 147, 159, 126, 113, 120, 146, 138, 126, 141, 132, 121, 131, 127, 122, 123, 109, 93, 129, 163, 156, 135, 137, 137, 134, 136, 140, 128, 121, 124, 124, 118, 116, 122, 126, 130, 108, 131, 132, 117, 115, 86, 73, 71, 105, 137, 158, 202, 188, 135, 115, 118, 121, 116, 121, 131, 128, 135, 121, 111, 120, 133, 121, 120, 101, 140, 108, 115, 141, 122, 105, 136, 145, 126, 127, 123, 113, 117, 117, 122, 121, 106, 74, 106, 109, 106, 106, 99, 91, 90, 103, 106, 111, 111, 115, 125, 130, 136, 140, 132, 120, 95, 94, 88, 87, 98, 124, 120, 126, 132, 123, 108, 104, 115, 115, 125, 114, 129, 127, 125, 127, 141, 133, 125, 120, 129, 140, 135, 122, 131, 125, 125, 127, 127, 135, 131, 126, 144, 149, 151, 140, 132, 125, 130, 130, 132, 129, 118, 111, 124, 129, 143, 145, 144, 137, 145, 144, 149, 149, 151, 149, 140, 158, 150, 156, 151, 158, 155, 154, 154, 157, 155, 149, 150, 154, 160, 153, 162, 163, 156, 157, 163, 158, 161, 165, 161, 168, 162, 156, 162, 167, 167, 163, 155, 162, 165, 163, 164, 159, 163, 169, 166, 157, 153, 160, 164, 164, 168, 161, 167, 156, 160, 156, 157, 158, 162, 153, 160, 156, 148, 166, 156, 152, 154, 153, 157, 152, 166, 156, 135, 142, 143, 136, 143, 134, 127, 143, 137, 150, 142, 143, 137, 123, 146, 139, 143, 127, 138, 159, 136, 136, 141, 136, 135, 141, 135, 132, 123, 134, 145, 130, 123, 131, 133, 121, 117, 148, 137, 130, 132, 128, 126, 119, 100, 97, 147, 156, 133, 135, 127, 146, 138, 131, 132, 132, 128, 128, 124, 122, 133, 133, 125, 131, 143, 143, 127, 127, 105, 81, 63, 99, 140, 122, 153, 180, 163, 132, 114, 116, 117, 116, 115, 122, 125, 125, 116, 126, 109, 147, 127, 126, 127, 122, 124, 129, 118, 90, 127, 141, 120, 120, 122, 118, 111, 124, 124, 131, 120, 104, 110, 108, 112, 101, 96, 94, 104, 100, 101, 111, 99, 107, 124, 135, 134, 127, 136, 130, 106, 101, 90, 90, 96, 112, 125, 117, 122, 124, 119, 115, 116, 116, 125, 124, 117, 124, 123, 119, 128, 129, 130, 126, 125, 141, 142, 127, 129, 124, 123, 123, 131, 133, 126, 131, 145, 140, 155, 137, 138, 118, 126, 136, 136, 124, 119, 114, 118, 127, 132, 140, 150, 145, 146, 148, 156, 147, 151, 148, 142, 152, 151, 154, 161, 157, 157, 155, 156, 157, 154, 149, 151, 150, 152, 154, 162, 157, 163, 160, 166, 156, 158, 155, 166, 158, 157, 159, 165, 167, 162, 157, 161, 158, 169, 161, 158, 156, 154, 171, 167, 162, 164, 169, 166, 167, 170, 164, 160, 162, 163, 156, 158, 163, 159, 146, 149, 154, 141, 163, 169, 154, 150, 155, 149, 157, 155, 144, 152, 145, 136, 139, 133, 135, 124, 141, 134, 139, 137, 147, 146, 130, 147, 146, 141, 122, 128, 153, 142, 136, 145, 137, 139, 133, 127, 139, 140, 127, 136, 138, 137, 133, 141, 122, 103, 130, 151, 132, 138, 125, 122, 119, 131, 110, 126, 130, 127, 128, 123, 133, 120, 124, 170, 128, 124, 125, 123, 126, 124, 133, 123, 135, 136, 144, 134, 137, 136, 103, 71, 91, 126, 127, 110, 147, 155, 162, 138, 122, 122, 105, 107, 119, 119, 119, 128, 124, 94, 147, 133, 131, 119, 136, 134, 132, 127, 118, 118, 122, 117, 124, 123, 124, 113, 117, 120, 131, 121, 108, 104, 100, 112, 106, 103, 102, 101, 98, 102, 115, 116, 114, 121, 110, 127, 129, 127, 120, 107, 114, 109, 100, 97, 108, 116, 114, 110, 115, 120, 116, 120, 103, 116, 121, 127, 125, 114, 120, 124, 130, 130, 125, 125, 130, 125, 123, 121, 115, 114, 116, 127, 126, 122, 116, 134, 140, 154, 140, 137, 124, 128, 129, 128, 131, 128, 124, 120, 132, 131, 132, 146, 152, 150, 147, 146, 145, 147, 149, 148, 157, 152, 143, 158, 160, 153, 159, 150, 153, 156, 150, 147, 135, 139, 156, 154, 152, 165, 157, 159, 159, 161, 159, 160, 158, 157, 164, 160, 168, 161, 166, 166, 164, 163, 159, 165, 161, 162, 164, 168, 170, 162, 165, 161, 167, 169, 159, 154, 158, 156, 154, 159, 156, 152, 146, 157, 155, 152, 149, 155, 143, 146, 160, 146, 145, 149, 149, 146, 142, 140, 131, 145, 131, 138, 138, 136, 148, 133, 144, 148, 142, 136, 145, 145, 138, 126, 150, 127, 135, 138, 141, 135, 136, 135, 132, 136, 128, 140, 137, 137, 114, 136, 141, 103, 121, 170, 126, 125, 130, 137, 126, 125, 118, 139, 130, 115, 130, 130, 130, 107, 107, 145, 132, 124, 126, 131, 116, 145, 135, 137, 142, 133, 133, 138, 135, 145, 128, 97, 89, 117, 116, 83, 106, 126, 145, 155, 136, 116, 127, 129, 121, 111, 120, 128, 124, 127, 128, 136, 132, 116, 133, 132, 128, 129, 130, 121, 134, 119, 122, 124, 118, 111, 121, 118, 129, 115, 111, 106, 97, 106, 106, 108, 102, 103, 107, 113, 109, 97, 144, 124, 116, 122, 123, 112, 103, 105, 116, 117, 107, 111, 117, 122, 120, 108, 107, 115, 120, 118, 120, 122, 119, 122, 125, 121, 123, 127, 129, 124, 121, 119, 117, 114, 126, 121, 113, 116, 114, 118, 127, 129, 132, 127, 119, 124, 123, 127, 131, 132, 138, 135, 132, 143, 138, 118, 119, 128, 137, 149, 146, 148, 151, 141, 139, 144, 146, 151, 148, 149, 151, 147, 153, 160, 159, 153, 152, 150, 155, 157, 149, 148, 157, 153, 156, 157, 153, 166, 149, 162, 161, 163, 158, 160, 156, 164, 167, 162, 159, 161, 156, 163, 159, 158, 165, 168, 164, 170, 169, 161, 169, 176, 163, 172, 158, 154, 156, 158, 153, 158, 153, 184, 145, 166, 153, 162, 148, 161, 154, 156, 156, 126, 130, 138, 136, 143, 136, 146, 128, 133, 144, 142, 145, 141, 148, 144, 138, 136, 141, 126, 135, 128, 150, 136, 137, 137, 139, 142, 145, 137, 141, 136, 130, 138, 116, 135, 144, 132, 115, 139, 161, 113, 118, 141, 120, 128, 121, 132, 130, 130, 103, 128, 165, 124, 107, 112, 133, 138, 123, 127, 131, 133, 131, 136, 137, 131, 142, 139, 142, 138, 141, 134, 141, 144, 136, 121, 110, 128, 115, 113, 99, 106, 114, 135, 141, 125, 128, 122, 127, 119, 124, 124, 130, 122, 123, 126, 125, 132, 127, 128, 128, 119, 125, 127, 127, 124, 108, 131, 117, 105, 108, 123, 124, 113, 102, 114, 109, 100, 98, 102, 95, 96, 126, 122, 96, 56, 146, 136, 119, 125, 121, 122, 108, 98, 110, 100, 104, 107, 119, 125, 117, 110, 109, 118, 116, 122, 119, 119, 121, 127, 124, 132, 128, 125, 133, 115, 119, 119, 103, 108, 128, 118, 116, 125, 109, 126, 127, 137, 138, 129, 125, 118, 114, 119, 122, 129, 135, 131, 132, 144, 150, 132, 121, 129, 132, 145, 141, 150, 145, 146, 146, 147, 151, 143, 151, 147, 152, 150, 159, 158, 153, 154, 154, 153, 151, 160, 161, 158, 154, 155, 157, 157, 155, 162, 157, 155, 154, 160, 168, 158, 159, 158, 161, 168, 164, 167, 164, 169, 162, 160, 163, 172, 170, 167, 165, 167, 171, 165, 163, 162, 160, 163, 154, 161, 160, 164, 122, 194, 155, 155, 159, 153, 153, 154, 160, 156, 153, 144, 137, 139, 148, 135, 127, 144, 140, 134, 143, 136, 144, 138, 140, 142, 141, 139, 136, 162, 131, 131, 142, 143, 138, 141, 138, 134, 145, 134, 145, 137, 141, 140, 137, 136, 135, 117, 87, 143, 182, 156, 133, 133, 123, 134, 124, 135, 132, 110, 74, 126, 181, 152, 93, 99, 124, 146, 131, 132, 112, 147, 131, 139, 144, 135, 139, 142, 141, 138, 144, 135, 139, 134, 128, 130, 111, 126, 115, 122, 115, 119, 126, 120, 126, 125, 129, 125, 123, 135, 111, 123, 132, 132, 128, 129, 121, 135, 132, 129, 118, 121, 123, 119, 120, 116, 116, 116, 125, 125, 132, 127, 110, 105, 96, 102, 91, 93, 98, 94, 92, 93, 131, 147, 120, 90, 103, 94, 117, 116, 111, 119, 122, 104, 99, 100, 95, 94, 121, 124, 112, 115, 112, 114, 117, 112, 119, 118, 124, 121, 128, 126, 126, 135, 141, 128, 124, 123, 115, 118, 109, 112, 119, 129, 121, 131, 133, 135, 134, 125, 121, 112, 121, 125, 124, 131, 130, 124, 124, 139, 139, 129, 130, 116, 128, 150, 149, 146, 148, 146, 143, 146, 151, 149, 156, 147, 139, 151, 155, 160, 146, 150, 152, 148, 157, 155, 162, 159, 156, 157, 158, 157, 157, 157, 158, 165, 156, 158, 165, 164, 171, 165, 162, 165, 164, 167, 162, 162, 163, 162, 164, 172, 165, 168, 164, 166, 169, 161, 164, 168, 155, 152, 157, 156, 160, 166, 155, 152, 161, 153, 162, 158, 159, 161, 148, 152, 155, 163, 149, 159, 138, 145, 126, 143, 133, 134, 136, 144, 146, 139, 148, 144, 138, 142, 134, 138, 133, 134, 143, 133, 132, 144, 138, 139, 141, 130, 149, 140, 130, 133, 134, 136, 130, 107, 87, 116, 170, 186, 168, 133, 123, 130, 129, 128, 140, 92, 62, 111, 177, 161, 106, 95, 122, 133, 123, 126, 114, 144, 139, 136, 137, 136, 133, 136, 141, 134, 136, 132, 152, 141, 132, 125, 127, 121, 118, 124, 121, 123, 137, 125, 127, 132, 119, 122, 124, 131, 118, 123, 122, 124, 125, 121, 124, 125, 118, 130, 122, 121, 122, 126, 105, 101, 115, 113, 121, 120, 138, 126, 109, 108, 103, 103, 90, 90, 98, 97, 78, 98, 109, 109, 119, 121, 111, 115, 123, 116, 116, 121, 119, 122, 107, 109, 105, 106, 120, 113, 117, 113, 108, 121, 114, 114, 110, 118, 114, 122, 120, 124, 123, 134, 135, 135, 128, 126, 118, 117, 109, 104, 116, 121, 124, 130, 132, 132, 131, 126, 123, 112, 117, 120, 126, 128, 125, 120, 116, 129, 130, 121, 137, 129, 137, 130, 150, 145, 147, 143, 147, 147, 143, 154, 151, 150, 151, 144, 154, 165, 128, 162, 149, 154, 157, 153, 159, 159, 159, 159, 149, 170, 169, 152, 159, 161, 166, 160, 159, 161, 163, 166, 163, 167, 164, 165, 166, 164, 161, 160, 163, 160, 169, 163, 168, 168, 165, 166, 165, 171, 159, 156, 156, 156, 162, 164, 150, 167, 165, 157, 140, 153, 154, 147, 161, 158, 148, 154, 155, 160, 142, 119, 120, 178, 132, 138, 141, 127, 143, 139, 145, 143, 142, 149, 144, 139, 139, 133, 158, 134, 114, 164, 135, 138, 138, 144, 134, 138, 141, 122, 137, 139, 119, 88, 93, 108, 156, 179, 197, 135, 119, 128, 119, 131, 125, 110, 46, 94, 140, 127, 106, 119, 127, 133, 123, 132, 115, 143, 132, 138, 139, 147, 137, 145, 141, 139, 144, 135, 140, 139, 129, 126, 126, 117, 116, 124, 116, 121, 130, 120, 121, 128, 120, 131, 135, 121, 125, 122, 130, 136, 133, 124, 134, 126, 112, 129, 117, 121, 109, 102, 133, 158, 119, 115, 126, 119, 126, 133, 130, 134, 117, 92, 66, 40, 82, 95, 84, 102, 110, 101, 109, 119, 121, 121, 115, 118, 117, 109, 116, 120, 119, 115, 107, 100, 113, 118, 119, 117, 103, 126, 107, 115, 107, 103, 106, 122, 125, 121, 116, 136, 138, 138, 133, 116, 121, 126, 114, 106, 117, 124, 126, 123, 133, 135, 129, 125, 126, 118, 112, 110, 128, 119, 120, 112, 107, 116, 122, 128, 127, 135, 138, 143, 139, 147, 144, 138, 148, 145, 147, 155, 149, 145, 146, 139, 148, 177, 149, 148, 153, 154, 156, 156, 158, 158, 147, 168, 149, 170, 155, 151, 160, 160, 163, 158, 156, 163, 157, 162, 166, 165, 165, 155, 167, 166, 162, 161, 155, 161, 165, 164, 165, 167, 164, 156, 156, 167, 161, 158, 159, 157, 149, 159, 145, 146, 141, 175, 173, 158, 167, 123, 160, 201, 170, 148, 154, 154, 137, 129, 130, 135, 145, 143, 113, 170, 133, 145, 130, 138, 141, 148, 134, 143, 132, 125, 132, 144, 116, 130, 139, 140, 129, 152, 141, 133, 132, 121, 138, 139, 104, 87, 100, 112, 141, 171, 194, 137, 123, 131, 132, 130, 137, 136, 109, 105, 113, 124, 130, 125, 123, 136, 120, 123, 122, 135, 134, 143, 132, 135, 146, 142, 144, 133, 135, 131, 138, 126, 126, 125, 120, 114, 120, 118, 112, 133, 127, 118, 132, 131, 126, 125, 133, 129, 123, 127, 131, 130, 132, 130, 134, 116, 110, 140, 152, 130, 98, 82, 127, 177, 160, 113, 118, 130, 129, 136, 135, 142, 130, 100, 80, 64, 78, 100, 109, 111, 106, 98, 98, 119, 113, 117, 115, 111, 103, 105, 113, 115, 112, 120, 108, 115, 115, 108, 115, 123, 114, 113, 109, 107, 103, 103, 116, 125, 128, 124, 121, 131, 130, 143, 132, 126, 125, 113, 112, 123, 118, 120, 125, 123, 123, 131, 130, 129, 127, 129, 127, 127, 121, 119, 118, 104, 100, 106, 104, 125, 123, 140, 147, 139, 143, 143, 147, 136, 143, 141, 151, 150, 145, 146, 144, 146, 148, 155, 151, 152, 152, 154, 153, 156, 162, 151, 154, 159, 154, 158, 138, 165, 161, 152, 164, 159, 162, 162, 158, 168, 162, 156, 162, 154, 166, 157, 156, 159, 157, 156, 161, 156, 160, 161, 166, 153, 161, 156, 154, 153, 151, 144, 156, 152, 157, 113, 121, 185, 193, 161, 160, 106, 144, 191, 178, 150, 156, 154, 149, 132, 125, 131, 141, 146, 72, 177, 124, 153, 138, 139, 148, 138, 138, 141, 136, 137, 140, 137, 126, 126, 141, 143, 135, 133, 140, 134, 135, 135, 134, 138, 93, 91, 96, 112, 130, 149, 154, 126, 120, 130, 130, 125, 129, 118, 135, 139, 129, 129, 131, 126, 126, 129, 130, 125, 119, 131, 139, 138, 142, 140, 143, 143, 142, 135, 132, 139, 112, 119, 127, 131, 117, 102, 109, 105, 105, 116, 121, 123, 120, 126, 125, 120, 127, 117, 122, 131, 131, 135, 130, 130, 124, 87, 83, 126, 161, 145, 109, 77, 126, 154, 143, 119, 121, 128, 126, 126, 136, 143, 123, 100, 90, 87, 84, 97, 104, 120, 116, 107, 102, 110, 122, 114, 101, 109, 123, 122, 111, 115, 112, 116, 107, 114, 100, 112, 105, 105, 97, 111, 111, 107, 104, 110, 133, 126, 126, 121, 121, 135, 138, 141, 136, 129, 120, 106, 95, 110, 115, 115, 114, 121, 117, 127, 126, 130, 122, 117, 126, 132, 120, 122, 113, 104, 77, 102, 105, 118, 110, 139, 153, 134, 142, 147, 146, 138, 142, 143, 154, 144, 153, 149, 143, 151, 151, 152, 147, 151, 150, 155, 153, 149, 166, 152, 166, 156, 134, 178, 150, 151, 158, 158, 163, 162, 160, 161, 158, 162, 157, 155, 158, 161, 155, 150, 151, 158, 152, 151, 150, 156, 153, 158, 149, 155, 148, 144, 147, 149, 146, 132, 163, 148, 145, 126, 126, 172, 151, 175, 163, 126, 143, 179, 163, 149, 157, 155, 128, 141, 136, 129, 124, 140, 134, 129, 136, 126, 144, 147, 142, 143, 147, 140, 124, 141, 136, 141, 135, 131, 128, 142, 123, 150, 131, 132, 133, 129, 133, 136, 112, 104, 98, 105, 114, 134, 124, 113, 136, 125, 138, 134, 124, 104, 128, 134, 121, 139, 128, 103, 131, 141, 135, 126, 121, 124, 135, 139, 141, 142, 143, 135, 130, 142, 139, 139, 115, 128, 136, 119, 129, 120, 111, 103, 114, 114, 107, 114, 126, 120, 129, 128, 127, 107, 120, 128, 129, 130, 135, 133, 127, 98, 68, 116, 135, 123, 125, 103, 108, 129, 125, 107, 114, 117, 122, 127, 122, 128, 129, 102, 93, 102, 94, 96, 106, 115, 115, 115, 101, 109, 113, 105, 72, 89, 126, 138, 122, 108, 112, 100, 96, 109, 103, 102, 95, 101, 98, 102, 116, 110, 116, 108, 117, 120, 104, 120, 125, 141, 155, 147, 143, 128, 126, 113, 106, 95, 100, 103, 102, 112, 114, 121, 121, 122, 130, 134, 126, 143, 124, 127, 119, 108, 93, 100, 99, 111, 114, 125, 128, 132, 145, 143, 143, 146, 139, 142, 146, 146, 149, 153, 147, 159, 156, 155, 154, 151, 150, 150, 154, 148, 148, 143, 173, 164, 127, 164, 160, 151, 157, 159, 156, 158, 159, 160, 158, 156, 159, 149, 163, 159, 147, 148, 152, 152, 147, 152, 150, 144, 144, 146, 143, 144, 142, 145, 143, 141, 137, 135, 139, 136, 144, 130, 150, 149, 138, 144, 135, 157, 169, 161, 151, 154, 153, 151, 137, 144, 138, 134, 119, 134, 125, 128, 137, 135, 140, 136, 146, 144, 130, 136, 136, 142, 135, 141, 135, 122, 138, 146, 128, 135, 136, 141, 137, 143, 133, 129, 135, 134, 120, 117, 119, 119, 109, 109, 128, 132, 139, 135, 136, 127, 130, 122, 125, 121, 132, 125, 121, 130, 129, 132, 129, 123, 133, 132, 136, 131, 136, 136, 137, 132, 138, 139, 133, 121, 122, 118, 119, 122, 115, 115, 123, 120, 103, 106, 121, 118, 127, 133, 129, 127, 129, 134, 130, 125, 126, 125, 122, 100, 73, 101, 126, 117, 119, 119, 128, 130, 125, 113, 116, 115, 130, 120, 118, 127, 126, 101, 105, 116, 100, 103, 115, 117, 114, 114, 102, 115, 111, 114, 71, 92, 113, 125, 110, 82, 94, 104, 105, 102, 105, 105, 102, 105, 114, 102, 119, 116, 118, 114, 113, 116, 77, 121, 125, 152, 148, 139, 142, 140, 134, 117, 117, 108, 98, 97, 84, 87, 92, 104, 109, 110, 131, 141, 144, 142, 135, 133, 116, 116, 111, 105, 88, 107, 110, 122, 130, 126, 138, 137, 142, 140, 132, 137, 147, 136, 142, 145, 186, 180, 159, 155, 154, 155, 149, 153, 158, 153, 135, 142, 166, 159, 155, 159, 160, 155, 164, 160, 153, 165, 158, 155, 156, 145, 153, 150, 152, 151, 134, 158, 176, 153, 149, 150, 149, 134, 158, 137, 124, 135, 139, 134, 147, 135, 143, 140, 131, 132, 142, 121, 159, 154, 143, 142, 144, 160, 142, 177, 163, 146, 148, 158, 129, 136, 134, 130, 124, 129, 127, 125, 139, 140, 149, 124, 142, 142, 138, 146, 136, 126, 133, 145, 138, 130, 137, 135, 132, 135, 131, 133, 136, 138, 145, 131, 130, 134, 131, 133, 135, 122, 119, 112, 127, 137, 128, 124, 137, 131, 124, 125, 127, 100, 124, 117, 118, 114, 124, 127, 124, 122, 130, 131, 134, 134, 128, 138, 140, 133, 128, 135, 129, 135, 133, 128, 120, 119, 113, 118, 133, 124, 109, 103, 120, 124, 128, 126, 133, 121, 122, 127, 118, 123, 121, 123, 121, 125, 112, 110, 123, 130, 125, 121, 128, 121, 125, 115, 121, 118, 114, 112, 105, 119, 110, 93, 111, 105, 109, 110, 104, 117, 103, 101, 108, 116, 105, 112, 91, 93, 99, 89, 82, 64, 102, 94, 92, 108, 104, 108, 103, 109, 106, 107, 108, 113, 115, 116, 104, 100, 95, 102, 123, 146, 146, 138, 143, 137, 134, 132, 116, 108, 100, 102, 94, 91, 88, 76, 81, 91, 116, 132, 140, 139, 140, 139, 119, 122, 117, 108, 105, 108, 103, 122, 123, 137, 135, 134, 140, 142, 139, 138, 147, 132, 132, 144, 200, 169, 149, 154, 157, 157, 146, 147, 152, 159, 153, 149, 157, 144, 153, 159, 152, 154, 151, 157, 143, 164, 156, 151, 153, 148, 142, 138, 147, 143, 141, 152, 150, 155, 148, 149, 155, 119, 164, 128, 116, 127, 134, 132, 129, 125, 133, 134, 126, 129, 137, 116, 142, 137, 140, 138, 157, 149, 140, 171, 165, 151, 155, 155, 142, 127, 123, 135, 138, 154, 127, 119, 153, 146, 140, 122, 132, 133, 137, 145, 136, 135, 136, 141, 129, 135, 139, 123, 140, 131, 124, 135, 137, 135, 138, 129, 135, 129, 125, 137, 137, 126, 130, 108, 132, 136, 130, 127, 140, 127, 131, 126, 135, 129, 130, 114, 121, 110, 131, 132, 119, 137, 139, 132, 132, 116, 116, 146, 153, 142, 130, 115, 122, 141, 140, 130, 125, 127, 128, 116, 118, 123, 124, 119, 127, 121, 122, 128, 134, 126, 121, 106, 108, 122, 132, 127, 129, 129, 127, 119, 120, 120, 122, 130, 127, 120, 119, 129, 125, 114, 105, 105, 106, 100, 89, 87, 89, 91, 117, 111, 115, 122, 109, 108, 118, 113, 104, 112, 111, 103, 101, 97, 80, 90, 106, 103, 104, 104, 109, 99, 95, 106, 102, 106, 103, 110, 95, 116, 112, 107, 104, 120, 131, 139, 142, 143, 149, 137, 135, 133, 121, 115, 112, 103, 97, 96, 93, 76, 74, 84, 94, 97, 116, 126, 144, 135, 130, 123, 121, 112, 111, 110, 109, 135, 126, 128, 136, 130, 133, 142, 134, 133, 141, 145, 136, 146, 163, 150, 150, 149, 153, 159, 132, 170, 143, 153, 153, 148, 147, 152, 143, 151, 151, 155, 146, 142, 147, 146, 144, 148, 150, 144, 135, 141, 136, 140, 145, 149, 139, 143, 145, 143, 141, 158, 139, 135, 130, 125, 124, 128, 141, 134, 132, 127, 129, 140, 145, 134, 130, 117, 142, 143, 159, 156, 155, 152, 155, 157, 150, 153, 148, 150, 124, 110, 134, 167, 142, 127, 136, 151, 130, 134, 118, 140, 141, 132, 144, 131, 136, 135, 129, 137, 133, 127, 122, 127, 130, 140, 134, 137, 133, 136, 138, 133, 125, 140, 130, 123, 129, 118, 131, 134, 136, 140, 136, 133, 125, 128, 137, 121, 131, 105, 82, 89, 124, 129, 123, 128, 133, 143, 127, 106, 108, 149, 163, 145, 127, 115, 124, 128, 132, 125, 128, 129, 123, 120, 121, 123, 130, 125, 122, 114, 107, 130, 131, 133, 114, 121, 121, 128, 136, 128, 135, 124, 136, 143, 128, 125, 121, 122, 123, 119, 132, 146, 138, 106, 115, 111, 94, 93, 85, 89, 91, 85, 98, 103, 115, 115, 114, 114, 110, 109, 103, 103, 108, 113, 112, 111, 90, 95, 109, 104, 103, 118, 111, 107, 95, 103, 104, 102, 107, 106, 107, 104, 113, 111, 107, 114, 123, 128, 138, 142, 138, 134, 130, 137, 129, 121, 109, 107, 110, 104, 106, 97, 81, 83, 79, 81, 72, 104, 133, 134, 134, 125, 125, 112, 121, 110, 110, 139, 128, 122, 126, 123, 127, 134, 129, 128, 141, 146, 142, 144, 145, 148, 143, 139, 157, 153, 130, 167, 150, 156, 159, 151, 148, 153, 151, 151, 152, 144, 150, 137, 133, 145, 145, 143, 143, 138, 135, 137, 133, 136, 141, 134, 142, 142, 140, 141, 129, 144, 130, 138, 131, 132, 127, 131, 142, 144, 145, 141, 138, 141, 148, 141, 149, 144, 148, 140, 152, 155, 158, 150, 155, 151, 151, 159, 143, 131, 100, 128, 141, 155, 122, 138, 129, 137, 132, 135, 129, 136, 137, 119, 144, 137, 131, 136, 131, 145, 129, 139, 134, 124, 137, 129, 131, 131, 127, 135, 139, 129, 126, 126, 140, 123, 140, 128, 122, 140, 117, 145, 131, 126, 129, 133, 134, 128, 125, 114, 104, 116, 132, 124, 134, 131, 131, 134, 133, 99, 121, 130, 149, 135, 140, 137, 134, 123, 127, 128, 120, 126, 130, 125, 128, 130, 129, 128, 120, 119, 108, 136, 124, 124, 125, 123, 113, 125, 145, 125, 125, 120, 134, 147, 133, 134, 144, 139, 130, 123, 126, 155, 147, 139, 135, 122, 88, 81, 89, 82, 78, 82, 85, 96, 107, 89, 95, 113, 111, 99, 91, 97, 105, 107, 110, 107, 101, 90, 98, 93, 91, 111, 106, 101, 105, 101, 100, 108, 110, 112, 123, 116, 115, 109, 114, 114, 113, 122, 127, 138, 121, 124, 132, 126, 128, 123, 117, 122, 122, 113, 109, 102, 93, 92, 92, 89, 83, 95, 120, 123, 133, 132, 120, 111, 119, 127, 128, 132, 129, 125, 133, 125, 128, 123, 121, 127, 138, 144, 137, 135, 146, 156, 146, 140, 155, 155, 158, 144, 151, 150, 151, 161, 157, 150, 149, 151, 159, 145, 134, 143, 128, 152, 136, 145, 139, 139, 136, 140, 138, 141, 137, 145, 141, 137, 140, 137, 129, 125, 140, 133, 134, 124, 135, 143, 145, 149, 139, 148, 149, 147, 145, 155, 148, 142, 157, 154, 157, 151, 152, 160, 149, 142, 149, 151, 131, 120, 145, 153, 159, 132, 126, 133, 136, 134, 135, 145, 133, 137, 141, 138, 142, 135, 148, 118, 155, 130, 141, 139, 138, 122, 137, 131, 141, 114, 132, 141, 139, 134, 138, 120, 141, 113, 133, 136, 107, 137, 135, 132, 133, 130, 128, 125, 127, 130, 125, 104, 91, 118, 124, 126, 123, 133, 124, 135, 137, 124, 122, 131, 130, 132, 130, 133, 136, 132, 133, 130, 121, 120, 133, 130, 124, 117, 129, 130, 119, 112, 107, 126, 128, 125, 124, 127, 122, 116, 135, 128, 119, 108, 131, 129, 118, 133, 147, 139, 131, 133, 122, 150, 155, 142, 138, 114, 79, 68, 80, 81, 77, 77, 105, 107, 109, 109, 120, 111, 106, 105, 98, 97, 99, 101, 112, 110, 113, 95, 99, 94, 87, 87, 89, 100, 94, 88, 96, 91, 113, 107, 109, 114, 111, 108, 112, 110, 115, 114, 119, 128, 134, 126, 128, 123, 134, 126, 131, 121, 129, 122, 111, 107, 112, 105, 109, 105, 100, 101, 109, 102, 114, 114, 105, 107, 116, 123, 137, 134, 128, 127, 131, 134, 126, 117, 111, 129, 135, 140, 139, 138, 132, 157, 149, 138, 149, 155, 152, 144, 157, 158, 140, 163, 156, 152, 152, 151, 143, 142, 144, 147, 137, 147, 138, 140, 153, 142, 134, 136, 150, 136, 135, 141, 141, 137, 127, 133, 129, 139, 143, 142, 138, 138, 131, 146, 143, 147, 152, 150, 153, 160, 141, 168, 156, 149, 154, 154, 163, 145, 160, 158, 153, 141, 164, 149, 124, 118, 149, 146, 147, 133, 140, 134, 134, 144, 142, 127, 142, 147, 133, 144, 141, 147, 140, 124, 128, 145, 146, 132, 146, 132, 134, 135, 133, 124, 132, 137, 141, 130, 139, 117, 124, 137, 134, 126, 122, 108, 135, 144, 133, 130, 124, 137, 133, 136, 131, 96, 122, 120, 115, 121, 127, 138, 122, 138, 138, 134, 131, 138, 129, 128, 121, 134, 132, 121, 131, 133, 126, 126, 127, 133, 130, 122, 116, 128, 129, 115, 117, 115, 116, 134, 130, 122, 125, 126, 126, 122, 123, 115, 112, 117, 118, 118, 128, 131, 135, 132, 125, 143, 152, 144, 137, 108, 81, 65, 67, 67, 78, 89, 95, 113, 119, 115, 113, 112, 111, 111, 104, 104, 100, 104, 114, 112, 100, 85, 98, 102, 90, 102, 102, 97, 88, 93, 102, 100, 111, 112, 106, 106, 94, 95, 115, 115, 114, 113, 121, 117, 129, 132, 123, 125, 128, 130, 131, 124, 132, 128, 121, 117, 122, 123, 115, 111, 108, 123, 118, 112, 99, 100, 110, 94, 100, 111, 123, 135, 147, 139, 133, 131, 120, 111, 106, 120, 130, 139, 131, 136, 153, 145, 148, 141, 153, 143, 153, 145, 150, 152, 152, 151, 152, 152, 148, 149, 144, 146, 142, 145, 145, 140, 134, 146, 144, 139, 134, 138, 141, 134, 139, 131, 133, 140, 135, 132, 144, 145, 138, 155, 139, 136, 147, 151, 152, 151, 160, 151, 151, 161, 160, 156, 153, 155, 159, 152, 159, 138, 172, 155, 160, 149, 145, 147, 121, 120, 150, 154, 124, 132, 138, 142, 132, 141, 132, 139, 135, 138, 146, 142, 137, 134, 144, 133, 140, 136, 141, 137, 137, 134, 140, 138, 137, 138, 139, 145, 145, 139, 127, 140, 127, 130, 125, 130, 120, 96, 114, 146, 135, 123, 126, 133, 130, 130, 126, 113, 112, 114, 121, 123, 131, 126, 127, 137, 136, 132, 135, 134, 126, 131, 134, 133, 139, 120, 132, 134, 131, 125, 127, 137, 125, 119, 116, 116, 130, 129, 122, 110, 113, 123, 116, 116, 121, 121, 119, 123, 122, 137, 119, 122, 127, 126, 119, 127, 128, 133, 135, 142, 157, 144, 131, 102, 75, 58, 67, 62, 70, 82, 98, 109, 112, 107, 110, 121, 108, 111, 108, 109, 98, 85, 103, 116, 97, 87, 95, 107, 83, 80, 97, 101, 99, 97, 96, 100, 115, 108, 104, 113, 93, 93, 111, 111, 107, 113, 107, 107, 117, 119, 127, 122, 125, 126, 127, 123, 133, 126, 124, 131, 124, 130, 117, 105, 119, 128, 124, 120, 104, 105, 127, 117, 97, 102, 106, 121, 144, 142, 144, 134, 124, 122, 115, 119, 126, 134, 123, 132, 159, 152, 147, 146, 150, 147, 151, 152, 148, 153, 153, 149, 152, 153, 151, 154, 154, 147, 146, 148, 143, 142, 151, 147, 139, 142, 132, 139, 142, 137, 139, 137, 136, 140, 138, 131, 146, 143, 137, 151, 141, 149, 155, 155, 153, 158, 157, 157, 152, 160, 164, 159, 157, 168, 168, 157, 167, 157, 147, 156, 156, 155, 153, 151, 117, 132, 155, 163, 115, 134, 128, 141, 142, 126, 135, 137, 129, 153, 141, 143, 133, 142, 150, 141, 133, 126, 145, 140, 135, 137, 130, 140, 137, 151, 140, 136, 141, 141, 145, 139, 130, 130, 132, 129, 120, 119, 116, 123, 134, 139, 142, 136, 124, 131, 126, 118, 113, 120, 113, 123, 134, 135, 137, 123, 136, 131, 132, 124, 121, 132, 137, 131, 136, 123, 126, 135, 129, 126, 108, 120, 133, 129, 124, 111, 118, 134, 130, 118, 109, 118, 114, 126, 120, 126, 121, 116, 110, 133, 122, 116, 122, 125, 126, 123, 132, 145, 148, 146, 155, 151, 126, 93, 74, 56, 66, 62, 64, 69, 92, 93, 98, 95, 103, 120, 110, 106, 111, 107, 96, 79, 93, 89, 92, 121, 110, 104, 94, 67, 93, 107, 93, 105, 110, 108, 107, 108, 103, 107, 89, 100, 109, 107, 92, 104, 105, 113, 105, 116, 113, 120, 127, 124, 124, 124, 127, 116, 129, 124, 136, 128, 127, 121, 119, 129, 117, 115, 109, 108, 132, 128, 107, 97, 98, 111, 132, 150, 152, 148, 134, 130, 124, 118, 122, 120, 123, 131, 144, 143, 148, 143, 139, 157, 131, 165, 155, 146, 143, 146, 149, 163, 156, 149, 152, 148, 152, 151, 151, 143, 145, 151, 140, 140, 137, 129, 132, 132, 143, 143, 146, 148, 145, 135, 146, 155, 150, 154, 137, 169, 152, 156, 157, 159, 158, 154, 159, 156, 162, 162, 162, 163, 160, 159, 166, 163, 158, 165, 160, 153, 155, 160, 114, 140, 144, 141, 144, 130, 133, 142, 140, 124, 156, 136, 135, 140, 135, 142, 141, 150, 144, 138, 130, 127, 118, 139, 137, 132, 147, 144, 121, 150, 169, 142, 134, 133, 145, 131, 121, 131, 137, 112, 128, 131, 127, 126, 120, 127, 130, 125, 119, 126, 124, 111, 110, 120, 120, 129, 125, 133, 136, 124, 125, 128, 129, 129, 138, 130, 143, 135, 134, 120, 141, 139, 131, 124, 126, 126, 122, 121, 120, 109, 112, 131, 128, 116, 92, 90, 113, 120, 124, 127, 122, 110, 118, 116, 113, 125, 127, 124, 125, 117, 113, 185, 160, 157, 161, 157, 131, 91, 70, 49, 61, 43, 49, 65, 83, 97, 100, 103, 103, 109, 96, 98, 102, 99, 93, 92, 97, 75, 76, 109, 119, 101, 97, 95, 105, 106, 96, 98, 95, 103, 110, 102, 100, 101, 97, 105, 105, 102, 95, 102, 104, 111, 117, 113, 101, 118, 119, 114, 120, 123, 116, 118, 130, 123, 126, 120, 120, 123, 131, 138, 128, 119, 111, 123, 122, 120, 120, 104, 86, 94, 108, 130, 156, 168, 150, 135, 118, 114, 122, 117, 132, 140, 145, 144, 143, 147, 145, 147, 131, 146, 169, 165, 148, 149, 143, 146, 150, 148, 150, 151, 151, 151, 151, 147, 143, 137, 145, 148, 145, 131, 143, 128, 142, 145, 148, 147, 147, 152, 152, 151, 153, 159, 118, 184, 166, 164, 158, 159, 158, 163, 162, 158, 163, 157, 166, 162, 163, 166, 161, 166, 157, 159, 163, 162, 146, 151, 135, 155, 134, 138, 125, 134, 130, 142, 131, 148, 128, 145, 139, 147, 141, 152, 138, 143, 141, 141, 142, 120, 149, 144, 134, 140, 138, 144, 119, 140, 158, 135, 129, 136, 139, 140, 134, 132, 125, 121, 125, 129, 108, 122, 128, 124, 122, 120, 120, 124, 124, 124, 111, 107, 116, 127, 127, 123, 131, 124, 124, 116, 122, 131, 140, 131, 129, 137, 125, 130, 128, 137, 128, 126, 127, 131, 127, 122, 124, 123, 123, 127, 135, 120, 117, 112, 119, 127, 116, 117, 121, 113, 108, 121, 117, 123, 129, 120, 126, 115, 90, 160, 154, 160, 164, 177, 139, 96, 69, 52, 55, 40, 43, 61, 61, 81, 90, 94, 92, 111, 117, 104, 98, 97, 94, 95, 100, 104, 92, 89, 91, 91, 99, 97, 98, 105, 97, 108, 117, 109, 101, 100, 124, 111, 101, 102, 98, 98, 94, 102, 109, 111, 116, 115, 113, 113, 111, 93, 107, 114, 117, 116, 120, 97, 118, 124, 120, 131, 132, 137, 141, 122, 109, 124, 118, 121, 125, 111, 87, 80, 94, 124, 148, 162, 149, 135, 116, 113, 106, 121, 126, 130, 144, 154, 143, 140, 149, 146, 124, 130, 160, 184, 153, 138, 156, 152, 144, 136, 148, 146, 143, 144, 145, 149, 139, 143, 152, 148, 138, 133, 158, 152, 145, 143, 143, 154, 156, 144, 155, 132, 153, 172, 140, 168, 155, 167, 158, 160, 158, 160, 159, 158, 159, 158, 159, 162, 169, 161, 163, 156, 155, 161, 162, 164, 156, 141, 143, 134, 132, 145, 137, 141, 129, 148, 136, 132, 133, 145, 121, 137, 143, 144, 146, 145, 146, 144, 137, 134, 133, 156, 141, 144, 132, 131, 140, 139, 133, 143, 131, 135, 144, 137, 136, 134, 126, 124, 130, 125, 125, 120, 109, 125, 124, 135, 126, 106, 128, 146, 141, 117, 125, 130, 135, 127, 115, 76, 147, 113, 121, 129, 131, 134, 130, 129, 128, 128, 128, 123, 127, 129, 125, 125, 129, 135, 125, 119, 131, 113, 128, 125, 118, 118, 115, 115, 124, 128, 122, 105, 106, 117, 115, 116, 113, 123, 129, 127, 120, 135, 142, 147, 166, 173, 151, 111, 64, 56, 65, 42, 36, 50, 55, 72, 75, 98, 99, 96, 105, 102, 94, 94, 93, 95, 104, 105, 102, 99, 110, 87, 94, 94, 105, 103, 100, 107, 112, 108, 88, 98, 132, 154, 119, 89, 102, 104, 107, 100, 101, 107, 101, 119, 120, 115, 120, 108, 106, 113, 112, 110, 103, 89, 116, 116, 128, 127, 121, 136, 136, 140, 126, 132, 128, 118, 122, 121, 92, 76, 86, 123, 148, 158, 147, 120, 108, 108, 110, 120, 113, 115, 141, 158, 150, 140, 132, 139, 147, 129, 151, 179, 150, 107, 161, 176, 144, 147, 151, 153, 148, 144, 145, 145, 137, 141, 151, 150, 146, 143, 152, 157, 146, 139, 155, 150, 153, 151, 167, 149, 151, 170, 147, 166, 159, 158, 163, 168, 160, 159, 165, 168, 159, 165, 166, 150, 158, 165, 161, 159, 160, 158, 157, 158, 163, 151, 149, 146, 135, 135, 132, 139, 137, 137, 125, 133, 137, 134, 135, 123, 141, 137, 145, 149, 146, 137, 141, 139, 142, 141, 138, 142, 140, 127, 148, 136, 142, 135, 134, 146, 132, 142, 143, 156, 119, 135, 123, 137, 132, 130, 116, 132, 122, 130, 120, 113, 118, 144, 138, 123, 120, 124, 132, 125, 128, 98, 113, 114, 115, 128, 132, 132, 128, 131, 127, 133, 125, 118, 125, 133, 131, 134, 127, 121, 129, 135, 125, 126, 117, 118, 120, 118, 121, 121, 109, 130, 126, 111, 117, 113, 115, 124, 112, 138, 125, 123, 123, 127, 153, 156, 167, 184, 175, 138, 79, 59, 59, 46, 29, 25, 31, 61, 81, 89, 93, 89, 109, 101, 94, 95, 82, 85, 106, 103, 90, 86, 99, 104, 97, 97, 94, 97, 99, 107, 105, 89, 70, 90, 122, 140, 119, 99, 105, 99, 97, 99, 75, 77, 91, 108, 115, 120, 123, 113, 112, 113, 119, 102, 97, 117, 125, 121, 135, 135, 153, 134, 138, 140, 138, 136, 136, 129, 126, 121, 101, 82, 87, 120, 138, 147, 133, 113, 103, 102, 106, 105, 107, 114, 128, 154, 158, 141, 121, 132, 163, 143, 142, 158, 145, 125, 143, 152, 145, 148, 147, 146, 150, 146, 149, 156, 149, 149, 150, 157, 150, 149, 153, 152, 154, 153, 151, 156, 152, 151, 159, 146, 166, 159, 166, 159, 160, 158, 157, 164, 158, 167, 162, 158, 156, 168, 161, 156, 161, 160, 161, 155, 159, 160, 152, 160, 159, 155, 131, 147, 136, 131, 141, 133, 139, 132, 146, 135, 131, 135, 136, 133, 146, 140, 136, 139, 147, 142, 138, 146, 143, 149, 129, 147, 146, 129, 142, 149, 136, 131, 128, 151, 133, 117, 129, 146, 134, 137, 127, 133, 105, 126, 127, 130, 128, 131, 120, 114, 119, 135, 116, 123, 131, 122, 130, 135, 129, 124, 126, 131, 115, 130, 135, 135, 128, 128, 128, 131, 121, 120, 116, 122, 135, 133, 127, 91, 111, 134, 101, 108, 123, 118, 119, 122, 115, 121, 123, 114, 114, 111, 119, 116, 120, 120, 108, 122, 123, 125, 122, 115, 130, 141, 159, 180, 187, 161, 116, 82, 53, 48, 34, 17, 14, 43, 70, 84, 98, 96, 105, 95, 88, 81, 76, 84, 103, 106, 100, 94, 97, 107, 110, 98, 90, 92, 90, 99, 103, 93, 67, 87, 114, 124, 102, 93, 103, 99, 95, 83, 64, 52, 88, 106, 106, 121, 118, 109, 114, 115, 116, 87, 91, 117, 124, 133, 137, 122, 129, 133, 138, 140, 151, 138, 139, 140, 136, 127, 114, 98, 100, 113, 124, 130, 119, 118, 104, 97, 101, 99, 112, 113, 128, 143, 151, 140, 128, 129, 159, 143, 134, 144, 146, 147, 142, 150, 145, 148, 151, 151, 152, 142, 155, 151, 155, 158, 154, 158, 158, 159, 154, 155, 149, 156, 151, 153, 158, 167, 167, 140, 172, 157, 158, 165, 163, 154, 165, 151, 162, 159, 164, 168, 158, 158, 165, 161, 162, 164, 157, 162, 159, 158, 159, 166, 167, 149, 137, 141, 141, 140, 131, 143, 131, 128, 139, 134, 135, 129, 131, 156, 137, 136, 140, 131, 138, 138, 147, 134, 148, 149, 133, 137, 149, 137, 137, 146, 134, 128, 132, 150, 137, 135, 128, 125, 136, 133, 115, 134, 123, 113, 122, 120, 118, 134, 123, 117, 126, 119, 116, 117, 128, 131, 124, 124, 120, 129, 133, 131, 123, 132, 133, 133, 132, 124, 124, 141, 132, 115, 123, 129, 130, 128, 125, 125, 126, 125, 120, 118, 119, 111, 105, 118, 124, 116, 115, 127, 116, 115, 112, 115, 120, 107, 115, 114, 119, 116, 115, 112, 126, 137, 150, 173, 168, 165, 116, 102, 78, 54, 38, 27, 18, 37, 69, 88, 107, 106, 102, 103, 85, 78, 81, 82, 98, 99, 95, 97, 89, 102, 90, 91, 90, 108, 98, 93, 86, 100, 90, 89, 100, 109, 90, 88, 102, 98, 102, 77, 52, 56, 72, 107, 103, 117, 116, 114, 117, 123, 118, 115, 108, 109, 113, 129, 131, 124, 128, 127, 138, 134, 138, 132, 139, 133, 136, 127, 124, 121, 124, 124, 135, 133, 120, 123, 111, 103, 93, 106, 114, 116, 134, 143, 138, 143, 141, 142, 149, 131, 131, 145, 150, 142, 147, 149, 154, 150, 154, 158, 151, 146, 156, 152, 158, 158, 156, 156, 154, 162, 156, 152, 155, 157, 149, 151, 164, 161, 161, 161, 156, 167, 160, 170, 173, 168, 166, 163, 159, 158, 164, 165, 168, 155, 168, 166, 153, 169, 158, 158, 163, 165, 153, 161, 160, 156, 140, 150, 146, 140, 143, 147, 141, 138, 137, 127, 143, 130, 136, 139, 133, 137, 132, 143, 132, 137, 147, 136, 146, 139, 138, 142, 139, 141, 144, 137, 123, 141, 144, 144, 142, 137, 131, 135, 134, 137, 141, 119, 134, 129, 124, 109, 105, 130, 129, 114, 118, 127, 122, 119, 119, 120, 110, 120, 109, 104, 129, 132, 127, 135, 132, 129, 129, 114, 120, 145, 116, 128, 118, 132, 123, 129, 126, 129, 126, 124, 126, 111, 120, 121, 110, 121, 117, 109, 104, 121, 117, 128, 111, 105, 111, 108, 113, 103, 103, 113, 109, 134, 118, 125, 138, 157, 164, 157, 130, 106, 91, 67, 40, 37, 31, 51, 73, 93, 106, 105, 104, 100, 80, 47, 43, 55, 69, 92, 103, 99, 92, 98, 95, 90, 91, 97, 105, 91, 94, 99, 98, 101, 108, 106, 100, 91, 102, 101, 94, 82, 54, 49, 73, 102, 113, 115, 112, 110, 115, 124, 122, 136, 121, 111, 116, 116, 118, 120, 137, 130, 134, 122, 128, 136, 139, 138, 132, 124, 122, 130, 135, 129, 140, 127, 123, 124, 107, 107, 105, 108, 113, 128, 135, 141, 141, 144, 143, 146, 148, 144, 143, 150, 151, 142, 148, 146, 157, 155, 156, 154, 149, 158, 159, 148, 154, 145, 150, 161, 157, 157, 157, 154, 152, 156, 159, 163, 164, 162, 155, 159, 156, 162, 159, 166, 165, 168, 169, 164, 161, 159, 170, 165, 165, 164, 164, 163, 163, 165, 162, 165, 158, 159, 157, 138, 156, 157, 132, 133, 140, 143, 138, 143, 143, 136, 140, 133, 138, 139, 137, 141, 127, 135, 142, 144, 146, 137, 142, 127, 155, 135, 141, 145, 151, 143, 136, 146, 136, 136, 153, 141, 138, 134, 135, 138, 129, 136, 131, 117, 125, 124, 120, 121, 117, 120, 124, 123, 113, 101, 113, 122, 115, 128, 112, 129, 124, 121, 127, 128, 132, 128, 134, 132, 125, 127, 126, 130, 124, 130, 124, 129, 129, 130, 128, 123, 125, 126, 125, 109, 110, 119, 118, 119, 115, 105, 97, 114, 104, 119, 112, 112, 120, 110, 119, 113, 108, 116, 103, 108, 116, 122, 135, 150, 152, 149, 135, 120, 109, 86, 63, 59, 57, 65, 79, 104, 105, 103, 93, 87, 73, 41, 49, 49, 54, 86, 92, 99, 95, 86, 98, 86, 89, 74, 89, 95, 103, 96, 97, 100, 100, 107, 111, 96, 93, 113, 99, 90, 74, 76, 87, 98, 115, 114, 122, 104, 120, 131, 126, 141, 128, 114, 127, 124, 124, 121, 137, 125, 130, 128, 125, 144, 137, 141, 121, 124, 124, 139, 139, 137, 139, 133, 120, 119, 113, 117, 107, 116, 119, 135, 144, 143, 131, 146, 152, 147, 144, 142, 147, 149, 152, 146, 150, 145, 159, 155, 155, 153, 152, 154, 157, 147, 157, 148, 152, 158, 160, 156, 161, 158, 154, 165, 158, 163, 166, 160, 168, 164, 161, 162, 165, 161, 161, 175, 165, 159, 155, 162, 170, 159, 171, 162, 149, 153, 156, 160, 173, 164, 152, 162, 155, 163, 150, 158, 136, 145, 132, 151, 142, 139, 137, 148, 143, 132, 131, 139, 130, 130, 126, 117, 134, 126, 150, 137, 133, 137, 133, 148, 149, 136, 136, 139, 140, 141, 131, 135, 147, 135, 153, 139, 136, 129, 138, 137, 128, 130, 122, 116, 101, 153, 121, 111, 129, 124, 109, 100, 93, 112, 110, 109, 115, 134, 104, 83, 122, 117, 124, 123, 133, 126, 115, 136, 128, 130, 125, 127, 123, 130, 119, 125, 126, 114, 124, 119, 125, 112, 111, 120, 117, 112, 118, 100, 109, 108, 112, 111, 114, 113, 118, 109, 114, 112, 108, 107, 118, 114, 111, 123, 130, 128, 129, 130, 127, 133, 118, 100, 87, 75, 73, 79, 97, 109, 114, 103, 100, 90, 73, 57, 53, 48, 53, 71, 87, 107, 86, 78, 91, 89, 86, 79, 84, 94, 94, 98, 92, 89, 103, 98, 113, 101, 96, 106, 103, 102, 104, 98, 93, 102, 112, 117, 120, 102, 114, 129, 133, 144, 132, 131, 139, 126, 129, 126, 125, 121, 125, 126, 129, 138, 131, 133, 128, 129, 130, 135, 142, 139, 137, 124, 117, 123, 123, 122, 115, 115, 119, 140, 141, 144, 143, 146, 136, 159, 140, 144, 146, 149, 149, 148, 150, 147, 153, 161, 149, 146, 154, 153, 151, 154, 164, 153, 150, 154, 158, 153, 161, 159, 160, 157, 164, 159, 153, 156, 163, 168, 167, 162, 163, 168, 155, 175, 164, 161, 162, 174, 165, 160, 164, 168, 146, 154, 159, 171, 159, 167, 157, 158, 155, 161, 152, 160, 148, 140, 143, 138, 143, 131, 141, 139, 139, 132, 133, 136, 125, 90, 165, 112, 143, 126, 133, 131, 134, 124, 130, 134, 124, 146, 168, 124, 132, 138, 132, 128, 129, 149, 139, 137, 147, 133, 115, 130, 122, 142, 118, 121, 87, 131, 116, 119, 129, 122, 120, 98, 91, 104, 124, 119, 120, 131, 118, 105, 106, 124, 125, 131, 118, 125, 123, 127, 122, 128, 127, 122, 120, 121, 124, 124, 128, 122, 119, 117, 118, 119, 111, 111, 113, 110, 111, 115, 107, 97, 113, 115, 118, 129, 115, 122, 103, 104, 108, 108, 107, 113, 106, 120, 130, 124, 119, 114, 110, 115, 132, 109, 105, 101, 96, 103, 99, 112, 122, 112, 104, 96, 69, 55, 46, 39, 66, 70, 88, 87, 86, 67, 85, 83, 81, 70, 87, 94, 91, 91, 94, 94, 109, 99, 95, 103, 104, 111, 101, 105, 104, 99, 106, 105, 113, 119, 117, 107, 108, 118, 127, 130, 127, 121, 145, 135, 132, 136, 133, 137, 122, 119, 130, 132, 124, 115, 127, 142, 129, 121, 138, 142, 132, 132, 125, 122, 127, 126, 120, 121, 130, 141, 138, 140, 150, 147, 141, 156, 149, 153, 143, 147, 147, 151, 149, 149, 151, 155, 152, 152, 166, 161, 150, 155, 155, 152, 156, 156, 154, 160, 161, 154, 159, 160, 172, 157, 167, 154, 167, 167, 158, 175, 167, 163, 162, 169, 161, 158, 162, 166, 161, 165, 171, 159, 158, 159, 169, 164, 167, 158, 149, 148, 165, 161, 153, 162, 140, 146, 136, 140, 135, 141, 141, 133, 138, 137, 137, 139, 61, 90, 204, 103, 116, 129, 136, 126, 142, 133, 125, 144, 108, 136, 178, 131, 136, 123, 137, 130, 137, 123, 147, 141, 135, 135, 130, 132, 138, 119, 131, 120, 115, 108, 132, 117, 116, 121, 120, 122, 107, 114, 125, 111, 118, 126, 120, 115, 104, 120, 118, 126, 123, 124, 131, 129, 121, 126, 122, 123, 118, 125, 131, 127, 123, 119, 121, 112, 116, 106, 109, 110, 110, 120, 108, 100, 117, 115, 116, 111, 109, 119, 114, 116, 107, 99, 101, 108, 126, 122, 107, 116, 127, 133, 114, 107, 110, 109, 110, 92, 110, 100, 105, 100, 99, 98, 123, 126, 102, 102, 61, 46, 44, 56, 62, 72, 83, 88, 95, 84, 86, 112, 93, 81, 92, 98, 96, 93, 83, 96, 98, 98, 94, 108, 105, 98, 96, 97, 103, 99, 101, 105, 111, 115, 118, 121, 111, 111, 114, 114, 114, 118, 134, 141, 133, 134, 130, 128, 123, 121, 128, 138, 127, 110, 126, 142, 132, 134, 139, 138, 127, 129, 129, 118, 128, 126, 116, 138, 136, 140, 139, 140, 151, 137, 153, 148, 151, 153, 144, 152, 156, 148, 155, 147, 145, 155, 156, 156, 197, 160, 155, 160, 149, 159, 155, 156, 166, 159, 161, 158, 144, 182, 171, 167, 161, 168, 169, 157, 165, 169, 164, 163, 168, 167, 166, 156, 158, 175, 156, 173, 168, 165, 169, 159, 158, 164, 162, 158, 160, 151, 172, 162, 152, 150, 132, 137, 127, 126, 137, 134, 142, 139, 139, 134, 141, 134, 48, 53, 162, 109, 129, 127, 135, 127, 129, 141, 121, 160, 132, 132, 133, 127, 135, 126, 131, 138, 133, 139, 140, 126, 139, 132, 132, 126, 132, 127, 127, 128, 115, 108, 123, 115, 117, 112, 117, 121, 123, 110, 95, 124, 124, 127, 130, 109, 113, 101, 116, 126, 114, 125, 131, 122, 127, 121, 118, 121, 116, 118, 120, 115, 110, 116, 118, 103, 115, 103, 96, 94, 95, 114, 113, 107, 110, 115, 110, 118, 118, 115, 108, 113, 108, 107, 109, 94, 141, 135, 115, 105, 122, 120, 117, 104, 109, 104, 114, 100, 105, 103, 105, 97, 92, 97, 111, 131, 98, 89, 71, 42, 42, 56, 68, 69, 88, 88, 93, 98, 97, 107, 99, 91, 97, 91, 72, 85, 82, 99, 99, 104, 107, 108, 98, 100, 100, 102, 101, 111, 99, 108, 109, 113, 124, 126, 125, 124, 118, 121, 109, 114, 129, 132, 134, 125, 129, 126, 125, 123, 138, 141, 135, 121, 126, 128, 130, 134, 135, 125, 124, 134, 127, 125, 132, 130, 125, 140, 141, 138, 138, 135, 145, 134, 151, 146, 144, 147, 141, 147, 152, 140, 159, 148, 144, 160, 157, 153, 172, 151, 154, 161, 150, 158, 155, 162, 160, 163, 157, 162, 156, 161, 163, 170, 158, 165, 165, 164, 159, 166, 168, 162, 171, 163, 162, 167, 161, 166, 154, 174, 168, 131, 177, 168, 161, 162, 164, 159, 164, 151, 170, 159, 168, 153, 121, 165, 188, 136, 137, 139, 147, 142, 141, 135, 105, 155, 127, 111, 107, 134, 118, 111, 137, 144, 134, 132, 128, 124, 136, 138, 138, 140, 134, 135, 135, 130, 138, 141, 142, 139, 135, 136, 129, 134, 133, 129, 128, 128, 121, 122, 118, 118, 126, 122, 108, 124, 118, 126, 121, 121, 126, 125, 118, 116, 102, 106, 135, 146, 124, 124, 111, 123, 123, 111, 119, 122, 113, 120, 112, 119, 106, 113, 116, 101, 107, 97, 81, 92, 103, 113, 122, 113, 110, 110, 120, 117, 112, 105, 110, 109, 103, 87, 106, 91, 116, 127, 113, 114, 107, 117, 108, 114, 102, 93, 121, 106, 102, 104, 111, 102, 94, 104, 113, 132, 113, 92, 80, 54, 48, 54, 68, 72, 74, 98, 101, 100, 104, 99, 102, 96, 98, 98, 88, 91, 90, 103, 105, 103, 105, 100, 93, 106, 102, 104, 101, 109, 106, 103, 110, 111, 123, 128, 126, 120, 122, 125, 122, 116, 130, 122, 127, 123, 119, 115, 116, 113, 123, 133, 138, 131, 133, 132, 129, 127, 130, 129, 120, 131, 123, 134, 135, 137, 140, 142, 142, 140, 137, 141, 147, 142, 142, 151, 147, 147, 148, 150, 147, 155, 149, 152, 149, 155, 158, 162, 159, 151, 160, 163, 155, 154, 158, 158, 157, 166, 159, 166, 164, 164, 163, 168, 167, 164, 165, 166, 148, 159, 165, 169, 168, 169, 160, 169, 161, 168, 169, 166, 164, 163, 165, 164, 169, 172, 168, 168, 163, 169, 170, 159, 164, 157, 119, 156, 185, 159, 133, 136, 154, 146, 138, 127, 123, 136, 131, 119, 124, 132, 128, 110, 130, 121, 148, 125, 127, 128, 132, 140, 136, 139, 133, 132, 148, 130, 161, 135, 134, 130, 141, 143, 130, 134, 136, 126, 119, 134, 134, 124, 118, 127, 102, 139, 136, 109, 112, 119, 109, 120, 125, 126, 110, 115, 99, 102, 121, 125, 120, 126, 124, 118, 117, 113, 122, 113, 102, 123, 116, 104, 99, 109, 108, 105, 100, 100, 108, 108, 105, 108, 109, 124, 113, 117, 116, 119, 105, 83, 116, 123, 101, 89, 102, 104, 110, 109, 118, 115, 112, 112, 117, 116, 110, 103, 105, 103, 109, 108, 115, 96, 86, 105, 113, 144, 115, 86, 75, 58, 53, 60, 69, 72, 77, 95, 103, 96, 85, 84, 99, 102, 103, 105, 89, 88, 105, 90, 96, 104, 106, 102, 105, 107, 101, 103, 107, 100, 118, 121, 116, 113, 123, 131, 127, 124, 111, 119, 121, 126, 135, 133, 128, 122, 124, 106, 100, 105, 118, 129, 138, 129, 134, 138, 126, 139, 130, 123, 129, 137, 133, 137, 136, 137, 134, 139, 131, 139, 131, 133, 143, 144, 139, 143, 142, 150, 149, 151, 147, 142, 175, 147, 151, 152, 156, 153, 158, 150, 156, 162, 158, 157, 155, 162, 166, 156, 165, 164, 159, 165, 165, 169, 164, 161, 164, 161, 157, 165, 163, 158, 164, 162, 159, 169, 161, 171, 170, 166, 162, 162, 162, 165, 160, 168, 162, 164, 159, 161, 167, 158, 163, 151, 119, 154, 170, 144, 136, 137, 136, 139, 135, 129, 139, 134, 108, 147, 126, 132, 126, 120, 126, 124, 124, 118, 125, 130, 136, 134, 137, 138, 132, 133, 130, 107, 152, 151, 133, 133, 133, 137, 131, 142, 140, 131, 111, 144, 138, 123, 118, 122, 73, 132, 167, 123, 111, 117, 115, 121, 130, 109, 114, 115, 102, 101, 111, 124, 111, 121, 122, 123, 119, 117, 121, 109, 85, 111, 134, 112, 88, 100, 110, 100, 89, 102, 105, 105, 105, 109, 105, 109, 126, 118, 120, 114, 98, 101, 112, 118, 110, 108, 106, 112, 106, 126, 113, 117, 106, 114, 113, 110, 121, 113, 102, 100, 113, 109, 114, 110, 96, 108, 118, 145, 136, 100, 80, 59, 60, 56, 66, 70, 73, 99, 95, 107, 92, 98, 94, 96, 96, 100, 103, 95, 96, 98, 93, 101, 106, 107, 104, 105, 109, 113, 107, 93, 108, 109, 116, 115, 111, 127, 128, 127, 118, 116, 114, 126, 143, 138, 132, 124, 118, 116, 96, 115, 123, 124, 128, 125, 124, 133, 132, 130, 130, 125, 131, 140, 138, 138, 133, 139, 139, 139, 134, 134, 134, 135, 145, 139, 137, 144, 147, 143, 144, 148, 147, 127, 164, 153, 146, 150, 150, 154, 158, 157, 155, 155, 158, 156, 153, 162, 163, 155, 167, 164, 161, 164, 169, 165, 164, 163, 160, 166, 158, 165, 168, 156, 162, 166, 161, 165, 165, 172, 165, 161, 166, 165, 158, 166, 161, 165, 169, 164, 161, 160, 153, 180, 165, 163, 100, 143, 150, 130, 137, 143, 144, 138, 119, 136, 151, 130, 106, 141, 127, 119, 134, 120, 137, 121, 133, 117, 125, 127, 130, 132, 141, 141, 133, 134, 142, 120, 130, 136, 137, 136, 134, 139, 129, 136, 140, 133, 117, 128, 127, 109, 110, 141, 106, 113, 127, 121, 125, 122, 86, 112, 161, 119, 116, 119, 114, 104, 104, 120, 118, 100, 107, 111, 116, 110, 112, 105, 84, 106, 122, 107, 101, 113, 114, 104, 108, 107, 98, 134, 107, 109, 118, 117, 114, 127, 128, 111, 107, 114, 118, 113, 109, 97, 98, 104, 91, 114, 111, 116, 104, 115, 112, 109, 122, 118, 114, 103, 114, 115, 116, 114, 108, 110, 133, 149, 135, 110, 76, 55, 49, 51, 61, 67, 73, 99, 102, 109, 109, 91, 89, 103, 98, 99, 110, 93, 76, 65, 81, 102, 100, 107, 103, 101, 100, 118, 102, 98, 102, 108, 108, 115, 115, 112, 130, 113, 110, 118, 126, 127, 134, 129, 132, 121, 118, 118, 112, 121, 123, 113, 124, 127, 119, 120, 123, 132, 130, 122, 139, 144, 142, 128, 131, 135, 139, 137, 144, 134, 126, 132, 136, 150, 136, 141, 149, 143, 145, 150, 145, 144, 147, 147, 146, 152, 146, 150, 157, 152, 152, 162, 156, 152, 157, 158, 164, 151, 160, 159, 158, 162, 170, 162, 159, 159, 162, 166, 160, 151, 162, 163, 160, 159, 163, 161, 168, 162, 172, 162, 163, 168, 165, 167, 166, 167, 173, 165, 168, 158, 122, 191, 167, 165, 120, 145, 137, 140, 141, 143, 141, 133, 123, 123, 146, 132, 123, 132, 126, 129, 127, 138, 123, 125, 119, 129, 130, 130, 128, 117, 150, 142, 131, 141, 127, 134, 117, 110, 124, 127, 134, 136, 91, 148, 133, 138, 126, 121, 120, 106, 107, 130, 126, 126, 105, 115, 115, 121, 84, 106, 135, 111, 115, 114, 117, 119, 110, 100, 114, 96, 99, 108, 116, 112, 114, 111, 101, 98, 103, 94, 108, 115, 118, 120, 101, 108, 100, 130, 127, 113, 116, 119, 111, 101, 121, 119, 103, 108, 115, 108, 104, 100, 89, 90, 101, 104, 110, 106, 100, 114, 113, 112, 126, 124, 119, 116, 124, 125, 120, 121, 119, 116, 142, 153, 142, 106, 79, 57, 45, 49, 62, 68, 69, 91, 98, 92, 101, 82, 98, 99, 100, 104, 102, 87, 86, 64, 89, 102, 103, 95, 107, 106, 101, 112, 104, 103, 111, 113, 110, 114, 111, 119, 118, 113, 109, 118, 128, 130, 127, 132, 126, 125, 118, 119, 120, 122, 121, 113, 124, 125, 119, 127, 135, 129, 128, 130, 135, 139, 127, 136, 142, 135, 142, 138, 143, 140, 138, 130, 125, 128, 144, 144, 144, 146, 151, 147, 151, 149, 143, 148, 149, 166, 159, 155, 152, 157, 148, 157, 156, 158, 160, 160, 165, 164, 158, 154, 169, 161, 168, 163, 158, 172, 167, 168, 163, 156, 164, 165, 162, 159, 163, 162, 159, 163, 166, 160, 159, 169, 144, 184, 159, 168, 168, 167, 173, 168, 159, 158, 157, 161, 133, 136, 140, 136, 130, 141, 139, 139, 128, 141, 135, 137, 132, 117, 122, 122, 127, 123, 124, 123, 133, 126, 115, 119, 130, 109, 131, 147, 127, 131, 117, 126, 123, 115, 111, 125, 135, 131, 120, 132, 131, 132, 115, 131, 129, 92, 114, 121, 109, 123, 129, 103, 113, 126, 111, 100, 126, 102, 93, 116, 99, 114, 116, 102, 107, 99, 104, 106, 109, 111, 113, 115, 112, 111, 110, 102, 113, 112, 123, 124, 107, 108, 105, 120, 124, 125, 95, 94, 112, 106, 98, 115, 125, 110, 96, 117, 112, 100, 94, 88, 103, 112, 104, 105, 109, 110, 118, 120, 121, 122, 128, 129, 123, 126, 129, 120, 114, 122, 132, 151, 151, 125, 84, 59, 30, 32, 54, 65, 77, 84, 83, 101, 103, 103, 101, 103, 105, 100, 100, 102, 88, 93, 98, 92, 99, 96, 105, 80, 90, 100, 111, 109, 113, 108, 116, 113, 107, 114, 109, 112, 108, 114, 123, 131, 123, 124, 128, 126, 124, 116, 130, 130, 122, 117, 119, 123, 121, 133, 127, 129, 130, 135, 141, 134, 100, 141, 164, 129, 143, 147, 144, 138, 134, 137, 132, 127, 137, 145, 139, 151, 149, 144, 149, 151, 146, 152, 144, 157, 158, 154, 152, 159, 148, 155, 154, 157, 155, 154, 162, 161, 158, 155, 163, 160, 158, 159, 165, 166, 157, 164, 160, 154, 155, 159, 167, 158, 151, 164, 160, 161, 160, 163, 162, 167, 159, 169, 161, 169, 167, 163, 161, 165, 165, 160, 162, 159, 137, 138, 139, 141, 139, 135, 133, 133, 132, 131, 126, 138, 124, 129, 126, 129, 132, 124, 128, 131, 122, 122, 120, 117, 111, 122, 119, 133, 127, 123, 114, 114, 128, 122, 122, 110, 131, 120, 131, 133, 134, 129, 124, 118, 141, 115, 103, 131, 112, 110, 129, 117, 94, 131, 138, 107, 118, 120, 102, 108, 117, 118, 117, 109, 93, 107, 107, 99, 110, 116, 110, 111, 111, 101, 122, 116, 118, 114, 124, 123, 114, 112, 116, 128, 118, 119, 115, 104, 119, 118, 107, 99, 118, 111, 114, 106, 112, 98, 105, 102, 102, 108, 104, 98, 109, 113, 114, 115, 115, 123, 140, 129, 131, 125, 127, 127, 120, 126, 120, 134, 150, 143, 112, 75, 26, 7, 34, 63, 80, 79, 88, 101, 105, 94, 94, 100, 95, 98, 112, 110, 100, 96, 102, 102, 97, 96, 103, 81, 94, 110, 115, 100, 95, 101, 110, 113, 109, 112, 115, 110, 109, 101, 118, 124, 131, 124, 124, 129, 121, 110, 125, 126, 126, 118, 122, 113, 119, 121, 127, 135, 141, 135, 129, 127, 121, 128, 142, 132, 139, 139, 142, 145, 139, 127, 144, 129, 138, 145, 137, 145, 148, 146, 143, 158, 153, 152, 150, 153, 142, 156, 153, 150, 154, 156, 142, 152, 154, 142, 153, 153, 159, 156, 162, 160, 159, 162, 165, 164, 158, 159, 159, 159, 158, 156, 162, 161, 166, 160, 157, 156, 166, 169, 160, 160, 169, 158, 157, 162, 160, 162, 162, 167, 165, 165, 160, 163, 141, 134, 138, 137, 126, 147, 141, 132, 125, 132, 136, 137, 130, 129, 129, 122, 125, 122, 134, 109, 105, 119, 159, 180, 126, 107, 105, 119, 121, 125, 133, 127, 126, 130, 123, 130, 135, 135, 126, 129, 119, 124, 137, 139, 118, 128, 118, 121, 117, 113, 112, 114, 102, 131, 128, 113, 98, 107, 108, 115, 106, 115, 111, 108, 102, 118, 116, 112, 106, 103, 105, 113, 119, 106, 112, 119, 112, 114, 115, 114, 110, 112, 121, 113, 116, 116, 115, 115, 106, 120, 125, 110, 112, 118, 116, 111, 112, 105, 107, 106, 102, 100, 109, 104, 106, 105, 105, 115, 114, 121, 123, 125, 125, 128, 126, 123, 129, 123, 114, 127, 139, 146, 129, 87, 27, 12, 32, 64, 78, 85, 87, 94, 96, 78, 96, 106, 92, 97, 103, 101, 101, 103, 119, 93, 80, 104, 108, 112, 106, 105, 116, 106, 112, 109, 109, 116, 110, 121, 116, 114, 106, 102, 110, 120, 128, 123, 124, 134, 123, 119, 112, 121, 127, 128, 120, 122, 123, 121, 127, 131, 132, 139, 138, 109, 142, 151, 136, 134, 134, 138, 144, 146, 142, 142, 146, 134, 141, 141, 141, 142, 154, 141, 143, 154, 147, 151, 160, 154, 150, 150, 152, 154, 157, 148, 154, 156, 153, 148, 160, 150, 144, 181, 159, 157, 156, 151, 160, 165, 159, 153, 166, 160, 156, 157, 160, 144, 175, 160, 153, 158, 160, 160, 159, 160, 164, 158, 165, 166, 163, 166, 162, 162, 161, 156, 161, 159, 150, 132, 143, 139, 137, 136, 141, 138, 132, 141, 126, 135, 136, 127, 127, 129, 130, 128, 121, 70, 88, 127, 153, 188, 201, 113, 99, 136, 116, 112, 117, 124, 122, 121, 133, 135, 126, 145, 117, 129, 110, 117, 112, 129, 108, 106, 138, 119, 112, 131, 117, 110, 114, 124, 122, 115, 112, 102, 117, 108, 106, 111, 117, 111, 106, 117, 103, 92, 117, 107, 106, 106, 111, 103, 103, 121, 120, 116, 124, 126, 109, 123, 125, 118, 111, 110, 103, 109, 116, 119, 117, 113, 113, 106, 105, 113, 114, 115, 115, 110, 109, 105, 108, 104, 99, 103, 108, 113, 119, 117, 127, 131, 130, 128, 126, 123, 133, 124, 120, 117, 131, 142, 137, 102, 52, 46, 47, 58, 81, 90, 93, 95, 96, 97, 100, 102, 102, 106, 101, 91, 77, 93, 121, 115, 103, 100, 109, 108, 114, 99, 117, 116, 113, 111, 104, 115, 121, 118, 111, 112, 104, 101, 110, 115, 115, 122, 121, 126, 127, 114, 100, 138, 126, 121, 111, 123, 131, 121, 125, 131, 130, 133, 140, 124, 122, 148, 136, 135, 136, 138, 140, 139, 141, 147, 148, 137, 150, 138, 133, 143, 143, 140, 152, 151, 143, 146, 154, 150, 144, 152, 156, 148, 155, 148, 142, 163, 155, 156, 156, 153, 123, 191, 158, 165, 158, 153, 159, 158, 170, 154, 161, 154, 159, 156, 156, 158, 155, 150, 157, 159, 158, 156, 166, 157, 165, 173, 157, 165, 164, 162, 165, 170, 168, 161, 161, 155, 140, 138, 141, 140, 140, 137, 143, 132, 137, 132, 134, 126, 139, 121, 127, 141, 132, 128, 126, 58, 83, 113, 142, 168, 213, 134, 100, 117, 107, 112, 121, 121, 127, 120, 130, 124, 114, 135, 119, 128, 114, 136, 118, 129, 105, 103, 127, 132, 101, 114, 118, 111, 118, 125, 116, 121, 118, 111, 118, 112, 87, 104, 120, 120, 110, 108, 106, 109, 93, 102, 106, 109, 109, 112, 102, 113, 118, 117, 118, 122, 114, 129, 130, 124, 117, 121, 118, 102, 123, 121, 117, 122, 106, 111, 110, 116, 123, 118, 115, 105, 105, 104, 103, 93, 92, 91, 93, 109, 110, 116, 123, 125, 128, 127, 131, 126, 130, 128, 118, 114, 131, 143, 123, 96, 70, 53, 59, 62, 75, 85, 93, 100, 92, 102, 102, 105, 103, 101, 96, 113, 98, 93, 94, 101, 104, 110, 115, 110, 112, 113, 114, 112, 117, 114, 108, 120, 118, 112, 99, 90, 107, 104, 112, 110, 116, 114, 124, 120, 120, 119, 106, 123, 114, 121, 121, 126, 128, 135, 129, 130, 132, 128, 131, 137, 131, 132, 137, 144, 140, 135, 139, 130, 138, 143, 141, 145, 144, 138, 140, 150, 146, 130, 145, 145, 150, 149, 149, 150, 151, 145, 144, 155, 149, 158, 145, 156, 152, 157, 153, 160, 139, 158, 159, 157, 155, 161, 152, 149, 160, 159, 162, 157, 154, 152, 155, 152, 157, 157, 161, 159, 165, 159, 164, 172, 163, 166, 158, 165, 161, 167, 160, 161, 166, 163, 161, 152, 139, 136, 139, 136, 140, 130, 145, 122, 127, 123, 132, 127, 132, 135, 126, 135, 131, 138, 113, 48, 78, 117, 143, 160, 196, 104, 114, 120, 120, 115, 115, 118, 118, 122, 133, 129, 127, 120, 129, 108, 129, 133, 128, 121, 112, 117, 124, 137, 125, 115, 118, 111, 105, 115, 111, 117, 116, 111, 115, 105, 101, 99, 104, 118, 105, 114, 119, 115, 111, 111, 99, 108, 99, 109, 118, 118, 121, 118, 114, 121, 130, 118, 116, 120, 123, 122, 116, 123, 120, 116, 117, 129, 110, 121, 113, 115, 112, 116, 116, 112, 106, 100, 103, 89, 81, 86, 74, 92, 103, 117, 126, 128, 130, 131, 128, 125, 123, 126, 117, 113, 122, 128, 111, 91, 75, 88, 66, 56, 72, 80, 99, 105, 89, 94, 103, 110, 110, 96, 102, 102, 104, 98, 103, 117, 108, 107, 104, 108, 116, 107, 111, 110, 114, 118, 121, 116, 115, 106, 90, 77, 101, 105, 114, 106, 118, 116, 124, 123, 124, 130, 122, 115, 116, 119, 121, 121, 128, 130, 130, 132, 130, 128, 122, 130, 138, 125, 138, 130, 144, 132, 140, 136, 134, 140, 147, 140, 154, 149, 144, 141, 139, 138, 139, 141, 148, 150, 150, 150, 155, 155, 154, 148, 153, 155, 149, 156, 155, 155, 155, 162, 150, 155, 157, 159, 158, 157, 158, 152, 156, 157, 155, 159, 151, 144, 148, 148, 151, 158, 156, 160, 160, 163, 159, 162, 157, 157, 156, 161, 161, 157, 165, 156, 159, 159, 158, 146, 140, 137, 134, 137, 133, 137, 132, 112, 99, 128, 142, 128, 113, 132, 128, 128, 126, 130, 129, 80, 67, 119, 128, 168, 138, 101, 120, 109, 127, 117, 118, 113, 134, 125, 111, 137, 122, 105, 138, 111, 129, 128, 122, 131, 101, 123, 127, 123, 131, 118, 111, 117, 108, 118, 115, 114, 116, 116, 108, 102, 100, 109, 114, 121, 104, 115, 119, 114, 119, 116, 117, 119, 107, 110, 118, 119, 123, 115, 116, 107, 124, 109, 108, 118, 114, 109, 104, 120, 119, 113, 115, 118, 89, 107, 124, 111, 124, 114, 107, 108, 89, 96, 113, 99, 90, 84, 72, 76, 84, 98, 118, 118, 126, 128, 124, 123, 123, 120, 125, 120, 112, 98, 98, 93, 114, 126, 94, 77, 73, 84, 96, 104, 101, 92, 106, 112, 111, 107, 109, 107, 102, 92, 90, 122, 110, 105, 105, 108, 115, 108, 111, 112, 110, 112, 123, 109, 110, 102, 101, 86, 98, 117, 112, 112, 113, 117, 121, 128, 128, 130, 125, 114, 120, 122, 114, 124, 128, 126, 130, 126, 128, 128, 131, 139, 135, 135, 133, 132, 136, 142, 143, 140, 139, 142, 148, 143, 153, 149, 144, 141, 138, 139, 149, 138, 142, 141, 152, 150, 158, 149, 155, 151, 153, 147, 148, 160, 154, 151, 163, 157, 149, 155, 157, 154, 157, 158, 159, 157, 155, 156, 152, 152, 149, 158, 149, 137, 167, 154, 160, 162, 161, 159, 160, 155, 166, 157, 154, 161, 158, 157, 156, 154, 160, 156, 154, 142, 143, 138, 132, 136, 135, 135, 134, 134, 128, 129, 130, 132, 132, 126, 129, 131, 106, 129, 117, 114, 86, 97, 114, 127, 105, 118, 121, 120, 121, 126, 119, 125, 123, 115, 137, 126, 101, 133, 122, 119, 121, 125, 102, 129, 116, 125, 114, 118, 119, 133, 115, 115, 129, 111, 110, 111, 111, 110, 111, 112, 104, 122, 116, 111, 117, 110, 99, 111, 117, 117, 114, 116, 107, 109, 114, 118, 114, 123, 109, 119, 116, 111, 114, 129, 119, 108, 102, 120, 111, 123, 119, 115, 113, 113, 114, 111, 115, 108, 107, 105, 102, 108, 120, 110, 101, 89, 70, 86, 81, 94, 107, 109, 108, 115, 121, 112, 111, 113, 117, 113, 119, 77, 73, 80, 126, 128, 116, 90, 76, 83, 97, 103, 99, 103, 102, 101, 105, 109, 111, 107, 95, 87, 94, 102, 109, 104, 97, 88, 104, 114, 108, 97, 118, 117, 125, 113, 109, 104, 107, 96, 105, 123, 119, 114, 106, 114, 117, 116, 118, 127, 120, 110, 113, 125, 123, 124, 121, 125, 122, 112, 130, 133, 136, 135, 139, 140, 137, 128, 134, 139, 133, 137, 140, 139, 141, 143, 143, 143, 152, 132, 151, 144, 149, 144, 138, 143, 154, 149, 148, 157, 150, 153, 163, 150, 152, 149, 155, 149, 161, 159, 153, 148, 152, 151, 159, 157, 153, 157, 151, 154, 150, 145, 157, 152, 137, 129, 177, 151, 154, 153, 158, 160, 161, 159, 152, 155, 161, 155, 156, 153, 155, 150, 158, 145, 150, 142, 133, 136, 131, 133, 134, 129, 132, 136, 135, 129, 127, 139, 127, 125, 135, 119, 115, 134, 130, 131, 143, 122, 123, 118, 116, 104, 122, 121, 126, 115, 106, 125, 116, 115, 125, 118, 105, 115, 115, 107, 133, 123, 146, 118, 116, 142, 123, 117, 115, 115, 124, 110, 120, 112, 102, 115, 119, 104, 104, 125, 117, 116, 117, 115, 119, 115, 109, 107, 105, 119, 112, 108, 121, 115, 120, 122, 110, 115, 124, 124, 113, 106, 137, 125, 109, 114, 114, 116, 117, 116, 117, 118, 111, 101, 103, 115, 114, 105, 87, 109, 123, 118, 117, 114, 99, 96, 87, 81, 85, 91, 96, 100, 103, 102, 106, 107, 111, 110, 117, 112, 120, 75, 61, 68, 99, 104, 101, 98, 93, 88, 102, 97, 102, 103, 95, 106, 101, 105, 106, 105, 98, 85, 116, 103, 105, 88, 105, 101, 101, 116, 108, 102, 105, 110, 119, 117, 111, 115, 117, 107, 107, 115, 109, 112, 116, 109, 114, 117, 116, 126, 119, 111, 123, 119, 118, 125, 121, 129, 129, 127, 120, 130, 128, 133, 127, 127, 137, 132, 131, 138, 134, 136, 137, 137, 141, 144, 136, 143, 152, 137, 148, 144, 148, 142, 146, 143, 151, 147, 152, 153, 144, 147, 150, 153, 152, 150, 148, 133, 174, 169, 159, 153, 155, 156, 150, 147, 156, 150, 155, 149, 155, 143, 143, 153, 143, 125, 157, 148, 153, 155, 160, 153, 157, 156, 162, 151, 152, 151, 148, 146, 142, 148, 143, 131, 140, 140, 137, 140, 134, 121, 125, 134, 130, 134, 137, 124, 133, 130, 124, 124, 123, 127, 120, 115, 128, 130, 134, 122, 125, 116, 120, 110, 122, 120, 121, 124, 120, 131, 113, 117, 118, 113, 114, 137, 116, 122, 128, 112, 141, 121, 116, 135, 125, 122, 115, 100, 126, 123, 102, 118, 142, 99, 116, 115, 95, 111, 121, 117, 121, 117, 109, 127, 125, 118, 119, 118, 117, 110, 114, 109, 110, 130, 121, 115, 125, 122, 108, 109, 130, 132, 122, 113, 113, 114, 108, 109, 115, 114, 101, 130, 110, 114, 114, 110, 101, 103, 148, 131, 113, 110, 116, 104, 94, 74, 72, 71, 77, 95, 100, 98, 103, 104, 108, 115, 117, 119, 130, 96, 63, 73, 99, 103, 90, 92, 91, 86, 107, 99, 107, 109, 104, 99, 105, 101, 115, 116, 109, 95, 103, 109, 112, 100, 93, 97, 106, 113, 95, 93, 97, 109, 112, 110, 121, 115, 111, 107, 111, 110, 114, 110, 115, 102, 91, 113, 114, 119, 117, 114, 126, 129, 128, 147, 131, 121, 136, 121, 113, 128, 134, 133, 127, 133, 128, 129, 135, 137, 137, 139, 140, 140, 143, 142, 141, 145, 149, 142, 149, 150, 148, 147, 151, 150, 156, 151, 146, 144, 149, 150, 152, 149, 146, 149, 148, 135, 146, 168, 168, 152, 153, 153, 149, 145, 151, 143, 151, 142, 152, 144, 124, 144, 156, 135, 145, 144, 157, 152, 149, 157, 150, 158, 153, 146, 151, 154, 151, 149, 137, 140, 134, 131, 149, 136, 135, 137, 131, 118, 117, 143, 137, 121, 137, 134, 134, 131, 113, 129, 119, 123, 127, 120, 119, 130, 128, 110, 132, 119, 119, 113, 114, 117, 124, 128, 116, 125, 131, 118, 124, 114, 129, 126, 118, 128, 136, 123, 127, 131, 112, 115, 128, 127, 114, 104, 112, 128, 111, 86, 148, 119, 105, 123, 97, 107, 113, 106, 119, 131, 111, 113, 124, 111, 109, 119, 115, 124, 118, 117, 107, 110, 118, 117, 125, 124, 111, 112, 108, 103, 111, 113, 109, 113, 113, 117, 115, 117, 111, 118, 107, 123, 119, 114, 103, 83, 134, 137, 123, 104, 112, 106, 95, 75, 68, 62, 59, 88, 98, 87, 103, 107, 101, 105, 114, 118, 126, 110, 82, 75, 98, 90, 87, 84, 85, 92, 110, 105, 108, 118, 115, 98, 111, 95, 98, 110, 103, 106, 105, 105, 111, 105, 109, 102, 110, 109, 92, 79, 87, 107, 102, 101, 111, 105, 109, 107, 103, 118, 117, 111, 114, 102, 81, 109, 117, 114, 119, 120, 105, 123, 119, 149, 126, 126, 133, 125, 128, 130, 127, 125, 134, 123, 129, 133, 131, 137, 130, 137, 131, 139, 140, 146, 142, 142, 147, 144, 149, 144, 149, 152, 144, 152, 150, 149, 143, 146, 142, 143, 147, 148, 148, 135, 173, 146, 144, 151, 149, 153, 128, 155, 147, 148, 152, 143, 141, 130, 138, 142, 130, 134, 145, 132, 139, 135, 159, 149, 143, 146, 150, 154, 156, 152, 152, 159, 150, 143, 144, 140, 128, 125, 146, 145, 144, 140, 131, 133, 132, 131, 137, 132, 136, 130, 136, 130, 117, 123, 133, 117, 124, 115, 115, 118, 146, 135, 126, 128, 112, 130, 128, 121, 129, 110, 124, 119, 120, 126, 112, 128, 121, 131, 121, 127, 131, 118, 127, 122, 112, 132, 119, 118, 125, 114, 119, 118, 123, 101, 123, 114, 125, 109, 60, 93, 140, 108, 117, 103, 145, 118, 121, 107, 117, 108, 113, 123, 123, 118, 119, 111, 113, 120, 122, 118, 115, 120, 112, 106, 117, 117, 124, 109, 97, 113, 116, 109, 112, 115, 100, 112, 115, 102, 107, 112, 138, 138, 126, 127, 118, 106, 92, 78, 66, 55, 49, 71, 89, 91, 94, 98, 96, 100, 117, 123, 122, 123, 110, 88, 95, 92, 79, 81, 82, 94, 102, 102, 112, 105, 107, 104, 104, 101, 101, 103, 106, 95, 117, 111, 108, 100, 98, 107, 104, 99, 91, 81, 92, 112, 110, 104, 107, 112, 95, 106, 113, 109, 108, 112, 112, 113, 103, 111, 110, 110, 90, 85, 77, 107, 121, 118, 116, 125, 130, 124, 123, 133, 127, 128, 132, 136, 138, 139, 135, 132, 130, 126, 134, 138, 143, 141, 137, 142, 147, 131, 161, 148, 148, 150, 141, 149, 152, 152, 140, 145, 145, 148, 147, 155, 153, 125, 165, 143, 153, 153, 147, 150, 139, 140, 142, 138, 136, 145, 134, 135, 137, 142, 143, 139, 136, 130, 135, 134, 148, 149, 150, 152, 153, 158, 143, 153, 144, 150, 150, 146, 148, 139, 136, 120, 135, 134, 120, 148, 137, 133, 137, 137, 129, 120, 119, 128, 134, 123, 130, 129, 125, 129, 117, 128, 123, 102, 134, 118, 127, 131, 123, 118, 119, 112, 132, 122, 121, 120, 120, 130, 88, 152, 128, 124, 124, 130, 125, 133, 133, 113, 135, 124, 132, 122, 123, 121, 128, 128, 122, 126, 121, 107, 116, 118, 99, 104, 123, 110, 120, 106, 118, 111, 121, 113, 114, 115, 111, 118, 116, 119, 114, 111, 110, 118, 118, 115, 117, 121, 121, 120, 116, 120, 119, 110, 92, 109, 113, 119, 116, 122, 109, 121, 116, 78, 69, 125, 170, 140, 130, 140, 131, 113, 88, 83, 61, 59, 58, 66, 79, 70, 69, 95, 103, 109, 123, 121, 122, 126, 124, 90, 94, 101, 90, 76, 79, 93, 106, 101, 95, 106, 103, 112, 112, 108, 107, 103, 101, 111, 111, 110, 107, 95, 92, 95, 104, 100, 106, 98, 105, 115, 121, 111, 116, 117, 110, 112, 118, 94, 104, 101, 114, 117, 116, 120, 120, 105, 85, 76, 77, 103, 114, 114, 116, 116, 127, 123, 120, 132, 129, 127, 133, 133, 132, 135, 134, 133, 131, 135, 140, 140, 148, 140, 141, 144, 145, 138, 150, 153, 135, 137, 144, 151, 143, 152, 134, 139, 149, 148, 145, 149, 151, 141, 137, 137, 152, 150, 138, 165, 149, 138, 143, 140, 143, 139, 140, 132, 139, 136, 134, 133, 136, 129, 136, 141, 145, 145, 153, 150, 156, 142, 147, 147, 139, 143, 139, 136, 136, 130, 136, 138, 144, 129, 132, 132, 138, 130, 134, 132, 95, 123, 136, 118, 139, 127, 125, 131, 126, 127, 127, 127, 135, 120, 133, 112, 120, 130, 120, 113, 136, 116, 124, 120, 114, 132, 121, 121, 123, 110, 128, 127, 117, 120, 121, 146, 134, 118, 115, 125, 134, 127, 125, 129, 123, 128, 110, 130, 120, 116, 105, 126, 122, 110, 111, 107, 111, 121, 123, 103, 104, 76, 97, 116, 122, 121, 118, 108, 102, 99, 102, 114, 121, 119, 112, 117, 116, 121, 119, 121, 124, 120, 117, 116, 117, 115, 114, 110, 116, 122, 116, 73, 53, 108, 153, 153, 141, 146, 137, 115, 106, 90, 63, 67, 67, 68, 69, 62, 60, 71, 95, 117, 129, 124, 121, 122, 132, 98, 95, 107, 96, 84, 69, 92, 97, 110, 109, 116, 104, 107, 105, 108, 104, 105, 107, 105, 100, 105, 111, 99, 98, 102, 103, 114, 113, 107, 108, 120, 114, 116, 117, 114, 109, 112, 114, 116, 110, 108, 113, 117, 119, 118, 113, 110, 102, 105, 107, 116, 115, 122, 121, 117, 126, 130, 128, 124, 129, 130, 135, 130, 128, 123, 133, 130, 137, 137, 140, 141, 144, 137, 140, 149, 143, 145, 140, 150, 142, 148, 158, 150, 146, 148, 146, 144, 142, 148, 146, 139, 150, 143, 130, 150, 152, 141, 117, 156, 153, 134, 138, 140, 139, 136, 131, 140, 136, 135, 137, 143, 137, 138, 142, 145, 149, 147, 152, 139, 147, 142, 143, 132, 129, 169, 139, 144, 135, 126, 137, 152, 136, 131, 135, 137, 137, 136, 131, 128, 37, 99, 183, 110, 131, 129, 131, 123, 124, 127, 129, 126, 126, 126, 127, 125, 119, 125, 122, 103, 144, 124, 108, 119, 119, 135, 99, 117, 122, 118, 129, 121, 111, 147, 122, 131, 118, 120, 119, 112, 129, 136, 129, 131, 116, 114, 116, 120, 125, 118, 121, 118, 114, 121, 125, 109, 126, 119, 121, 110, 109, 109, 91, 92, 106, 128, 120, 114, 109, 103, 97, 110, 114, 120, 119, 116, 118, 114, 107, 119, 116, 121, 119, 113, 116, 118, 114, 109, 112, 124, 120, 76, 54, 97, 136, 146, 146, 138, 133, 120, 107, 90, 79, 68, 67, 68, 62, 56, 56, 66, 81, 112, 135, 135, 126, 115, 119, 105, 104, 108, 98, 89, 79, 94, 97, 88, 116, 141, 105, 98, 101, 102, 104, 100, 98, 103, 99, 109, 111, 101, 98, 104, 101, 111, 114, 120, 118, 108, 107, 101, 110, 107, 115, 115, 111, 114, 109, 116, 116, 121, 117, 113, 106, 113, 111, 110, 110, 124, 109, 112, 118, 136, 124, 137, 134, 127, 116, 122, 135, 131, 129, 121, 130, 124, 133, 132, 140, 141, 140, 140, 141, 140, 146, 137, 141, 140, 143, 148, 148, 152, 149, 147, 150, 140, 138, 139, 148, 147, 139, 151, 145, 138, 148, 148, 132, 146, 149, 148, 133, 142, 137, 139, 136, 131, 136, 132, 138, 142, 133, 142, 147, 146, 146, 148, 161, 141, 144, 140, 134, 150, 143, 153, 133, 143, 145, 137, 150, 139, 141, 135, 134, 131, 131, 144, 137, 136, 89, 72, 113, 116, 135, 120, 130, 120, 126, 133, 130, 124, 127, 127, 121, 129, 118, 126, 121, 113, 127, 116, 122, 117, 128, 129, 115, 118, 119, 111, 135, 128, 116, 131, 131, 127, 98, 130, 110, 141, 124, 136, 126, 126, 131, 119, 110, 114, 118, 123, 117, 117, 116, 111, 116, 115, 122, 116, 113, 120, 115, 119, 110, 109, 112, 125, 117, 119, 111, 103, 100, 106, 115, 115, 116, 102, 110, 119, 102, 116, 115, 129, 122, 124, 106, 122, 125, 117, 109, 114, 127, 107, 87, 96, 123, 133, 140, 138, 121, 118, 104, 89, 94, 75, 75, 64, 59, 47, 50, 56, 68, 100, 128, 130, 118, 115, 128, 117, 101, 111, 96, 90, 94, 98, 97, 88, 104, 136, 109, 105, 104, 103, 107, 106, 92, 99, 107, 100, 103, 115, 116, 102, 105, 104, 108, 91, 117, 137, 102, 95, 104, 99, 115, 108, 115, 110, 109, 108, 112, 118, 110, 119, 116, 116, 111, 113, 99, 111, 116, 111, 106, 136, 126, 129, 128, 129, 133, 127, 127, 133, 126, 130, 125, 136, 133, 134, 143, 143, 142, 140, 143, 135, 145, 137, 140, 144, 150, 155, 147, 148, 150, 146, 149, 139, 146, 145, 147, 142, 147, 141, 145, 145, 149, 143, 146, 132, 138, 152, 137, 135, 138, 133, 134, 126, 136, 136, 142, 138, 138, 145, 148, 141, 125, 143, 169, 149, 142, 141, 138, 137, 146, 144, 147, 146, 146, 143, 151, 145, 144, 124, 133, 143, 136, 135, 131, 131, 129, 119, 123, 131, 134, 120, 141, 138, 132, 127, 135, 142, 118, 125, 118, 127, 123, 119, 121, 128, 122, 125, 114, 122, 128, 128, 131, 127, 123, 122, 121, 136, 125, 135, 128, 128, 134, 130, 129, 135, 131, 124, 130, 125, 128, 126, 123, 122, 116, 127, 115, 88, 115, 122, 113, 116, 120, 120, 120, 119, 114, 117, 118, 110, 125, 132, 117, 119, 109, 104, 106, 105, 110, 118, 125, 117, 112, 114, 119, 116, 118, 121, 114, 122, 128, 99, 123, 140, 110, 123, 125, 117, 105, 86, 121, 128, 148, 149, 113, 111, 105, 101, 100, 97, 80, 75, 65, 49, 40, 46, 62, 89, 117, 116, 114, 113, 113, 107, 105, 104, 110, 106, 97, 101, 93, 86, 101, 127, 119, 110, 97, 100, 105, 100, 101, 96, 93, 91, 104, 121, 137, 96, 95, 102, 115, 100, 86, 131, 110, 105, 104, 117, 118, 119, 113, 106, 102, 109, 114, 117, 115, 120, 117, 110, 115, 110, 107, 108, 108, 114, 110, 129, 122, 127, 129, 121, 133, 131, 126, 135, 132, 121, 118, 130, 139, 138, 136, 137, 134, 139, 138, 145, 134, 134, 142, 144, 144, 150, 150, 147, 147, 142, 147, 147, 147, 139, 145, 141, 146, 118, 159, 143, 147, 143, 145, 128, 135, 154, 143, 138, 145, 138, 131, 129, 131, 136, 138, 134, 139, 141, 144, 146, 141, 142, 155, 137, 137, 134, 147, 144, 138, 147, 147, 146, 150, 150, 148, 154, 147, 137, 139, 135, 137, 139, 129, 135, 135, 133, 139, 143, 137, 120, 116, 172, 134, 118, 131, 135, 118, 125, 126, 116, 132, 125, 119, 127, 126, 129, 125, 133, 107, 145, 135, 116, 127, 126, 134, 108, 121, 125, 130, 127, 134, 132, 140, 131, 132, 133, 129, 124, 127, 127, 128, 124, 127, 113, 115, 113, 108, 110, 107, 103, 102, 112, 115, 119, 119, 120, 115, 107, 113, 124, 115, 118, 109, 111, 107, 105, 105, 112, 123, 115, 108, 103, 119, 124, 116, 123, 121, 125, 125, 109, 111, 133, 119, 120, 111, 115, 114, 105, 107, 109, 134, 143, 123, 114, 103, 108, 107, 113, 94, 74, 75, 59, 32, 19, 61, 90, 104, 99, 110, 104, 109, 116, 109, 101, 125, 112, 101, 102, 103, 98, 102, 97, 118, 101, 117, 104, 97, 125, 102, 108, 104, 85, 93, 116, 118, 94, 103, 105, 108, 115, 117, 123, 109, 124, 117, 117, 118, 115, 114, 110, 104, 112, 89, 105, 119, 114, 118, 116, 112, 115, 108, 108, 110, 121, 119, 120, 111, 125, 125, 117, 124, 133, 122, 128, 131, 118, 125, 130, 140, 133, 133, 137, 134, 142, 143, 137, 147, 138, 139, 141, 135, 144, 147, 147, 144, 143, 152, 148, 143, 142, 141, 138, 144, 134, 136, 138, 139, 135, 145, 113, 137, 159, 146, 116, 157, 130, 131, 134, 127, 131, 138, 138, 133, 141, 141, 150, 146, 156, 148, 147, 141, 150, 136, 149, 128, 147, 145, 146, 146, 148, 141, 142, 150, 144, 137, 136, 138, 130, 142, 139, 131, 124, 138, 132, 133, 138, 114, 147, 132, 127, 139, 132, 129, 131, 125, 125, 116, 120, 113, 113, 118, 114, 117, 126, 86, 131, 157, 104, 129, 112, 124, 121, 118, 125, 156, 129, 129, 130, 126, 124, 127, 130, 89, 149, 118, 128, 125, 122, 122, 122, 116, 108, 101, 112, 102, 117, 106, 115, 110, 104, 120, 120, 118, 112, 122, 125, 117, 121, 114, 120, 117, 114, 100, 111, 118, 118, 117, 113, 113, 116, 110, 119, 123, 126, 125, 126, 129, 120, 114, 127, 109, 104, 113, 119, 120, 115, 125, 124, 113, 109, 106, 110, 129, 108, 96, 85, 80, 76, 57, 54, 69, 82, 96, 103, 98, 80, 100, 109, 103, 97, 112, 110, 103, 98, 98, 106, 109, 91, 97, 70, 101, 106, 113, 131, 118, 107, 113, 103, 96, 114, 103, 90, 104, 110, 117, 110, 111, 118, 116, 122, 116, 113, 112, 116, 118, 105, 127, 113, 103, 117, 117, 112, 121, 114, 109, 113, 114, 103, 116, 111, 126, 121, 127, 126, 117, 126, 120, 130, 130, 128, 119, 122, 128, 122, 131, 126, 135, 135, 138, 137, 137, 125, 141, 135, 144, 138, 142, 141, 146, 145, 149, 141, 142, 141, 141, 138, 142, 132, 135, 136, 141, 140, 141, 139, 148, 131, 135, 144, 139, 124, 147, 127, 128, 139, 129, 125, 132, 140, 142, 139, 151, 155, 152, 150, 152, 145, 139, 151, 141, 140, 147, 147, 143, 141, 150, 134, 145, 137, 156, 143, 128, 136, 133, 132, 139, 135, 136, 130, 132, 130, 135, 143, 113, 143, 131, 131, 139, 132, 115, 131, 125, 111, 122, 112, 108, 121, 105, 114, 105, 114, 122, 127, 97, 101, 119, 99, 108, 141, 111, 91, 141, 139, 128, 128, 130, 125, 123, 128, 109, 116, 136, 125, 126, 125, 118, 115, 112, 121, 114, 93, 109, 105, 93, 96, 121, 105, 114, 110, 111, 115, 117, 118, 117, 117, 114, 120, 121, 120, 110, 108, 125, 119, 109, 122, 119, 116, 122, 119, 126, 118, 122, 115, 124, 126, 120, 116, 114, 104, 112, 112, 121, 118, 128, 129, 106, 103, 93, 93, 137, 108, 95, 83, 78, 79, 65, 71, 70, 74, 82, 94, 87, 89, 97, 99, 113, 120, 108, 117, 108, 98, 102, 110, 114, 109, 95, 73, 84, 97, 112, 113, 102, 112, 111, 110, 103, 97, 85, 96, 96, 115, 118, 115, 114, 111, 114, 118, 109, 110, 104, 117, 110, 106, 110, 107, 117, 116, 115, 115, 113, 104, 114, 108, 115, 106, 113, 127, 128, 130, 145, 121, 112, 122, 128, 125, 129, 131, 126, 123, 126, 132, 134, 132, 136, 137, 130, 138, 135, 135, 133, 135, 139, 146, 144, 144, 152, 140, 147, 145, 145, 145, 140, 133, 140, 132, 135, 136, 141, 135, 140, 138, 141, 140, 139, 128, 133, 142, 125, 140, 130, 125, 137, 121, 145, 141, 135, 138, 151, 144, 144, 140, 149, 147, 142, 138, 151, 144, 151, 159, 149, 147, 145, 148, 140, 147, 158, 146, 131, 137, 139, 132, 134, 131, 134, 113, 132, 137, 133, 131, 117, 135, 137, 134, 139, 131, 134, 117, 128, 124, 115, 106, 117, 124, 115, 116, 99, 101, 124, 112, 107, 139, 115, 103, 99, 122, 117, 122, 116, 127, 125, 135, 148, 132, 135, 125, 129, 131, 124, 127, 125, 126, 131, 125, 120, 117, 119, 113, 110, 106, 73, 140, 121, 119, 120, 116, 112, 109, 113, 110, 104, 111, 118, 123, 118, 121, 122, 113, 124, 118, 111, 108, 113, 113, 117, 123, 122, 125, 124, 110, 116, 109, 109, 118, 110, 107, 124, 125, 120, 105, 115, 128, 105, 105, 97, 95, 100, 102, 102, 84, 79, 84, 73, 74, 79, 85, 74, 74, 85, 90, 108, 111, 111, 118, 113, 114, 105, 104, 84, 111, 119, 112, 88, 101, 112, 94, 100, 100, 94, 106, 111, 111, 112, 109, 97, 99, 95, 107, 112, 110, 105, 99, 112, 111, 96, 105, 115, 115, 108, 103, 103, 99, 116, 112, 108, 107, 108, 99, 115, 123, 118, 114, 117, 120, 120, 130, 143, 123, 110, 123, 129, 125, 131, 123, 134, 131, 128, 130, 130, 131, 128, 134, 133, 135, 126, 129, 137, 133, 139, 146, 138, 143, 141, 140, 142, 135, 143, 142, 145, 139, 146, 132, 141, 138, 135, 131, 136, 132, 140, 136, 138, 128, 135, 136, 122, 138, 133, 131, 126, 120, 141, 145, 145, 138, 145, 146, 145, 144, 146, 152, 140, 141, 145, 140, 145, 149, 145, 148, 146, 148, 149, 160, 154, 148, 130, 138, 137, 134, 137, 133, 123, 137, 137, 132, 130, 128, 135, 128, 124, 135, 135, 130, 142, 114, 137, 121, 123, 117, 118, 111, 126, 115, 109, 98, 121, 116, 129, 103, 109, 119, 118, 111, 118, 135, 121, 135, 138, 123, 120, 135, 125, 138, 126, 137, 128, 133, 130, 131, 129, 126, 112, 119, 110, 107, 127, 121, 106, 120, 118, 118, 114, 109, 116, 110, 118, 116, 116, 109, 117, 117, 112, 114, 125, 118, 124, 126, 122, 107, 114, 119, 116, 120, 120, 124, 117, 107, 118, 110, 117, 118, 113, 101, 116, 117, 128, 107, 110, 131, 138, 107, 102, 87, 74, 75, 104, 94, 64, 98, 89, 86, 94, 91, 74, 61, 74, 95, 109, 110, 112, 114, 103, 101, 95, 103, 103, 117, 121, 114, 86, 99, 138, 114, 98, 107, 112, 105, 103, 102, 119, 148, 142, 108, 109, 107, 113, 114, 111, 110, 105, 99, 109, 93, 111, 104, 120, 106, 108, 108, 111, 98, 108, 113, 107, 112, 112, 118, 116, 106, 117, 116, 120, 129, 144, 129, 114, 120, 137, 135, 134, 139, 124, 126, 126, 123, 133, 138, 117, 130, 131, 136, 134, 134, 133, 136, 141, 144, 140, 138, 143, 135, 133, 131, 143, 143, 145, 131, 141, 142, 129, 138, 130, 136, 134, 135, 133, 134, 139, 136, 136, 127, 127, 126, 131, 128, 132, 136, 133, 139, 149, 148, 136, 143, 148, 155, 146, 145, 139, 143, 143, 150, 146, 152, 149, 160, 151, 154, 154, 151, 154, 157, 133, 130, 136, 133, 145, 132, 118, 139, 132, 125, 125, 136, 131, 134, 128, 128, 135, 137, 136, 101, 142, 121, 117, 128, 112, 115, 99, 105, 115, 115, 120, 96, 131, 108, 118, 111, 123, 125, 132, 123, 134, 130, 130, 137, 134, 139, 132, 133, 131, 141, 127, 130, 124, 130, 128, 123, 125, 122, 118, 123, 117, 114, 119, 115, 114, 111, 97, 111, 105, 130, 121, 116, 117, 104, 108, 123, 119, 124, 123, 122, 118, 129, 126, 121, 113, 116, 113, 116, 105, 127, 109, 112, 109, 113, 112, 121, 115, 110, 111, 120, 121, 121, 118, 123, 123, 118, 97, 81, 66, 57, 85, 92, 72, 81, 93, 108, 95, 83, 72, 48, 45, 82, 114, 122, 107, 104, 109, 108, 106, 112, 114, 107, 113, 116, 94, 91, 108, 117, 108, 111, 109, 107, 102, 93, 119, 146, 163, 126, 109, 102, 104, 106, 106, 110, 106, 99, 111, 110, 115, 108, 110, 99, 129, 117, 109, 108, 102, 110, 111, 117, 112, 109, 112, 110, 113, 117, 121, 125, 137, 129, 105, 110, 123, 123, 122, 124, 120, 112, 126, 115, 120, 130, 128, 132, 130, 129, 136, 133, 134, 133, 140, 147, 141, 137, 149, 139, 136, 125, 134, 146, 147, 142, 143, 124, 143, 137, 134, 150, 133, 130, 132, 135, 138, 134, 134, 133, 119, 126, 123, 130, 129, 139, 136, 138, 138, 146, 145, 145, 152, 151, 149, 141, 150, 150, 151, 146, 144, 139, 150, 153, 151, 152, 159, 155, 159, 156, 132, 138, 129, 122, 130, 139, 128, 119, 120, 130, 135, 132, 139, 140, 134, 142, 122, 125, 130, 137, 124, 116, 108, 125, 117, 110, 91, 84, 83, 95, 117, 117, 112, 116, 120, 113, 121, 113, 129, 136, 131, 127, 123, 132, 128, 130, 124, 130, 103, 123, 133, 137, 121, 122, 111, 116, 120, 117, 110, 118, 140, 122, 117, 111, 138, 119, 117, 123, 66, 114, 129, 97, 102, 107, 103, 121, 113, 120, 127, 107, 92, 155, 112, 116, 118, 108, 111, 115, 111, 115, 111, 120, 107, 112, 119, 109, 107, 115, 115, 115, 113, 115, 129, 124, 124, 125, 102, 65, 38, 57, 76, 82, 80, 76, 72, 109, 115, 86, 73, 62, 66, 73, 94, 118, 97, 108, 110, 110, 112, 107, 107, 114, 106, 107, 112, 100, 110, 107, 113, 117, 104, 103, 97, 84, 115, 148, 141, 118, 110, 101, 106, 102, 108, 112, 106, 114, 118, 98, 113, 108, 109, 96, 109, 103, 108, 113, 111, 110, 105, 115, 105, 108, 110, 118, 118, 114, 112, 119, 131, 106, 116, 110, 121, 121, 131, 123, 118, 114, 118, 115, 129, 127, 129, 125, 127, 126, 127, 134, 127, 136, 145, 139, 143, 138, 144, 134, 139, 134, 130, 133, 142, 144, 129, 137, 136, 130, 135, 140, 161, 141, 131, 141, 139, 144, 138, 137, 125, 123, 123, 131, 128, 140, 140, 138, 133, 146, 143, 145, 147, 158, 150, 145, 157, 147, 149, 146, 148, 150, 150, 159, 149, 151, 164, 151, 154, 149, 126, 137, 128, 134, 137, 126, 129, 118, 126, 126, 140, 138, 135, 132, 121, 145, 131, 127, 121, 123, 118, 118, 110, 111, 109, 103, 98, 101, 108, 99, 110, 110, 113, 125, 121, 117, 126, 124, 103, 125, 128, 136, 122, 129, 139, 138, 135, 126, 110, 124, 133, 127, 132, 126, 119, 119, 122, 116, 113, 82, 136, 123, 125, 86, 131, 120, 117, 118, 121, 115, 115, 112, 101, 102, 112, 117, 118, 126, 114, 122, 86, 129, 113, 113, 117, 111, 103, 107, 103, 114, 112, 118, 106, 107, 108, 120, 114, 101, 99, 97, 105, 124, 125, 115, 113, 120, 111, 75, 39, 54, 87, 89, 86, 77, 61, 103, 135, 96, 78, 73, 77, 83, 86, 102, 97, 105, 113, 104, 112, 110, 100, 110, 110, 107, 112, 103, 106, 110, 111, 117, 107, 105, 108, 91, 109, 129, 125, 107, 100, 100, 110, 107, 105, 97, 106, 106, 113, 106, 109, 105, 110, 103, 104, 99, 106, 109, 102, 107, 104, 105, 107, 101, 112, 118, 115, 117, 118, 122, 127, 124, 121, 116, 129, 124, 143, 133, 114, 125, 123, 124, 122, 130, 134, 125, 126, 128, 122, 135, 126, 127, 144, 140, 142, 136, 138, 138, 135, 134, 137, 141, 139, 137, 133, 136, 139, 132, 138, 137, 142, 136, 127, 134, 136, 133, 136, 133, 122, 121, 125, 129, 128, 143, 134, 143, 139, 147, 148, 149, 141, 149, 145, 151, 151, 146, 148, 145, 149, 159, 153, 155, 166, 158, 163, 163, 155, 152, 132, 143, 126, 130, 132, 142, 134, 131, 136, 134, 132, 140, 132, 126, 134, 131, 133, 134, 121, 125, 116, 122, 114, 121, 117, 101, 107, 108, 111, 110, 109, 122, 115, 114, 120, 120, 111, 135, 131, 135, 135, 133, 101, 125, 133, 130, 144, 141, 122, 132, 135, 133, 128, 116, 131, 125, 123, 117, 119, 119, 123, 107, 126, 114, 109, 112, 112, 109, 119, 113, 102, 117, 102, 103, 116, 115, 118, 111, 113, 127, 128, 114, 115, 117, 108, 108, 101, 110, 107, 101, 105, 104, 101, 109, 121, 112, 113, 109, 100, 86, 89, 113, 128, 122, 111, 106, 124, 96, 73, 68, 81, 95, 103, 85, 60, 83, 99, 80, 78, 72, 79, 80, 86, 96, 101, 105, 109, 111, 111, 104, 104, 107, 107, 115, 114, 113, 101, 102, 119, 118, 115, 107, 86, 114, 109, 122, 106, 98, 95, 110, 105, 105, 115, 102, 109, 108, 105, 110, 91, 92, 102, 113, 108, 114, 108, 98, 100, 99, 94, 97, 109, 104, 110, 103, 106, 121, 114, 121, 116, 123, 122, 113, 119, 119, 124, 120, 124, 120, 124, 121, 119, 130, 121, 121, 126, 123, 118, 124, 126, 129, 136, 135, 132, 142, 135, 137, 135, 129, 137, 138, 138, 137, 140, 131, 132, 135, 138, 132, 134, 136, 129, 137, 134, 126, 126, 119, 126, 121, 126, 134, 138, 139, 144, 141, 149, 150, 148, 152, 153, 147, 143, 153, 147, 145, 150, 148, 156, 156, 157, 164, 155, 151, 164, 160, 159, 165, 136, 132, 131, 128, 133, 127, 132, 134, 125, 136, 129, 130, 133, 128, 129, 138, 127, 130, 119, 116, 108, 107, 127, 119, 102, 114, 109, 115, 106, 108, 110, 120, 114, 122, 125, 117, 101, 111, 110, 133, 130, 134, 85, 136, 136, 131, 140, 137, 124, 144, 132, 136, 121, 128, 126, 128, 127, 124, 119, 127, 124, 114, 121, 120, 120, 122, 110, 114, 124, 109, 84, 113, 121, 107, 122, 112, 115, 116, 118, 126, 110, 104, 116, 109, 107, 108, 107, 102, 100, 99, 103, 94, 109, 112, 115, 118, 115, 107, 112, 84, 67, 100, 113, 119, 121, 120, 118, 109, 84, 69, 71, 95, 113, 105, 90, 83, 83, 81, 75, 78, 75, 75, 82, 87, 104, 108, 110, 114, 105, 109, 111, 110, 100, 114, 110, 101, 113, 105, 105, 129, 112, 112, 106, 122, 117, 120, 113, 114, 100, 96, 101, 102, 113, 96, 99, 107, 104, 102, 105, 104, 96, 117, 103, 108, 103, 100, 100, 91, 82, 98, 104, 101, 111, 110, 105, 118, 113, 113, 107, 114, 113, 118, 121, 125, 119, 118, 120, 120, 114, 128, 118, 115, 116, 117, 116, 119, 119, 126, 126, 129, 129, 136, 128, 137, 132, 128, 134, 138, 143, 136, 128, 129, 134, 138, 136, 135, 140, 132, 129, 127, 134, 129, 127, 126, 113, 111, 114, 124, 134, 133, 136, 137, 146, 146, 150, 149, 150, 146, 145, 158, 149, 155, 153, 149, 145, 152, 152, 160, 158, 158, 164, 160, 155, 154, 160, 157, 130, 138, 133, 128, 137, 128, 130, 130, 130, 141, 134, 131, 132, 129, 139, 137, 125, 134, 119, 116, 114, 118, 119, 110, 106, 112, 102, 106, 114, 106, 109, 111, 116, 111, 123, 118, 88, 161, 119, 127, 137, 135, 129, 137, 136, 128, 144, 132, 137, 135, 139, 140, 126, 128, 130, 129, 114, 121, 127, 115, 117, 113, 116, 116, 126, 131, 121, 122, 118, 117, 93, 102, 112, 116, 88, 141, 121, 113, 115, 115, 100, 97, 100, 105, 97, 112, 94, 97, 105, 107, 110, 104, 104, 111, 110, 107, 116, 119, 111, 103, 95, 97, 108, 103, 106, 133, 145, 121, 102, 78, 62, 79, 101, 102, 111, 112, 92, 69, 81, 95, 65, 66, 76, 87, 107, 117, 112, 115, 108, 110, 118, 105, 90, 110, 109, 102, 114, 109, 104, 113, 108, 113, 112, 110, 107, 117, 122, 120, 101, 97, 96, 107, 109, 98, 91, 91, 98, 95, 104, 95, 92, 118, 105, 98, 87, 107, 103, 100, 92, 86, 100, 107, 98, 127, 110, 115, 113, 111, 111, 105, 121, 126, 121, 129, 120, 112, 100, 124, 125, 117, 112, 113, 114, 116, 119, 117, 125, 126, 125, 128, 134, 122, 126, 127, 121, 120, 135, 140, 139, 141, 131, 127, 135, 135, 133, 134, 135, 137, 133, 132, 135, 122, 116, 135, 113, 105, 114, 119, 127, 139, 140, 140, 146, 145, 150, 150, 156, 149, 154, 149, 150, 147, 143, 150, 154, 154, 162, 160, 161, 161, 161, 165, 166, 159, 163, 164, 137, 128, 129, 135, 135, 119, 125, 120, 136, 137, 137, 132, 130, 128, 125, 135, 127, 125, 120, 129, 131, 116, 118, 109, 101, 130, 105, 88, 114, 109, 123, 124, 119, 110, 126, 107, 99, 130, 126, 138, 126, 134, 138, 131, 146, 137, 135, 132, 137, 133, 129, 136, 129, 124, 138, 119, 130, 117, 107, 129, 103, 118, 119, 128, 124, 121, 121, 109, 121, 120, 108, 108, 115, 116, 88, 110, 115, 115, 113, 113, 107, 102, 94, 107, 102, 107, 103, 109, 108, 120, 108, 107, 116, 118, 110, 99, 118, 120, 124, 104, 84, 106, 98, 89, 97, 130, 143, 129, 110, 95, 82, 75, 84, 87, 100, 126, 117, 80, 73, 76, 51, 67, 79, 82, 107, 112, 124, 112, 108, 109, 111, 125, 109, 111, 114, 110, 114, 107, 103, 108, 117, 114, 109, 116, 105, 106, 125, 111, 113, 99, 99, 91, 90, 103, 123, 100, 96, 108, 105, 102, 111, 99, 103, 104, 101, 118, 97, 86, 92, 101, 94, 101, 79, 111, 108, 118, 112, 101, 119, 105, 112, 119, 125, 119, 118, 90, 96, 118, 124, 110, 103, 112, 104, 95, 124, 129, 126, 126, 123, 125, 129, 118, 129, 124, 91, 121, 131, 139, 134, 139, 129, 133, 134, 131, 137, 132, 137, 134, 131, 124, 134, 124, 105, 119, 109, 103, 112, 126, 123, 133, 145, 139, 144, 142, 134, 147, 163, 148, 150, 152, 149, 150, 149, 150, 154, 162, 157, 162, 165, 164, 162, 157, 146, 185, 160, 164, 133, 135, 133, 137, 134, 127, 133, 129, 134, 136, 129, 129, 128, 140, 124, 132, 129, 126, 126, 129, 119, 126, 122, 108, 110, 110, 101, 101, 110, 112, 120, 115, 101, 109, 100, 137, 95, 120, 117, 125, 124, 125, 138, 131, 145, 135, 136, 132, 130, 127, 124, 137, 134, 113, 131, 121, 121, 103, 105, 107, 126, 114, 123, 114, 91, 147, 110, 121, 109, 106, 108, 106, 115, 111, 100, 104, 107, 104, 110, 106, 108, 106, 107, 105, 112, 110, 107, 118, 112, 111, 112, 111, 114, 120, 109, 115, 121, 114, 105, 99, 87, 98, 94, 98, 110, 118, 122, 124, 105, 83, 76, 79, 80, 72, 103, 109, 102, 83, 80, 66, 55, 73, 81, 97, 107, 106, 117, 110, 111, 101, 93, 116, 137, 115, 102, 111, 105, 111, 109, 109, 107, 110, 118, 116, 105, 117, 115, 104, 110, 99, 94, 72, 57, 98, 135, 117, 92, 112, 97, 103, 119, 108, 97, 102, 102, 94, 103, 96, 84, 100, 100, 104, 89, 103, 100, 107, 107, 101, 106, 103, 105, 106, 118, 125, 119, 94, 97, 114, 96, 84, 99, 109, 107, 108, 123, 123, 117, 121, 114, 125, 126, 124, 134, 130, 117, 122, 135, 124, 136, 135, 134, 135, 140, 136, 134, 134, 133, 136, 128, 126, 134, 128, 103, 109, 106, 103, 106, 115, 127, 136, 139, 144, 142, 146, 145, 150, 157, 147, 151, 142, 156, 157, 156, 150, 140, 170, 159, 167, 158, 161, 150, 171, 146, 163, 166, 160, 147, 135, 136, 128, 148, 127, 137, 132, 129, 140, 129, 133, 120, 137, 127, 131, 132, 131, 124, 128, 129, 121, 118, 120, 118, 123, 117, 116, 126, 115, 119, 115, 127, 113, 108, 101, 123, 103, 125, 126, 142, 126, 135, 126, 141, 132, 129, 132, 137, 122, 126, 129, 131, 126, 130, 129, 128, 122, 113, 110, 116, 123, 129, 124, 69, 133, 114, 124, 113, 111, 115, 86, 117, 124, 102, 87, 106, 107, 107, 114, 106, 111, 114, 119, 112, 116, 111, 113, 116, 114, 113, 110, 117, 118, 108, 104, 114, 110, 108, 91, 97, 99, 103, 106, 107, 122, 117, 100, 97, 87, 73, 81, 77, 90, 108, 99, 92, 73, 65, 52, 60, 70, 79, 98, 106, 112, 122, 108, 108, 102, 90, 105, 125, 130, 114, 120, 104, 111, 101, 101, 113, 102, 107, 100, 95, 121, 107, 103, 106, 93, 107, 70, 47, 82, 121, 107, 96, 104, 96, 107, 108, 101, 100, 100, 106, 101, 96, 98, 95, 88, 104, 92, 97, 108, 111, 99, 98, 104, 104, 106, 102, 99, 109, 115, 118, 114, 97, 89, 82, 82, 75, 91, 108, 123, 124, 119, 113, 125, 119, 120, 131, 128, 126, 130, 130, 122, 124, 127, 136, 129, 132, 136, 131, 130, 134, 127, 139, 129, 128, 129, 116, 124, 109, 109, 110, 100, 103, 122, 133, 146, 138, 145, 149, 149, 147, 154, 152, 149, 143, 152, 178, 164, 153, 159, 149, 156, 158, 167, 164, 162, 161, 171, 164, 156, 167, 170, 142, 140, 139, 92, 142, 133, 128, 128, 118, 136, 135, 127, 132, 140, 133, 133, 128, 120, 140, 133, 121, 125, 118, 129, 128, 108, 125, 127, 124, 124, 118, 117, 106, 140, 122, 116, 122, 120, 117, 139, 130, 120, 140, 128, 138, 131, 136, 133, 128, 125, 127, 130, 125, 124, 128, 128, 131, 133, 119, 115, 115, 126, 124, 127, 129, 126, 116, 118, 112, 107, 104, 88, 108, 110, 104, 102, 111, 90, 106, 110, 110, 98, 99, 113, 110, 119, 113, 115, 116, 109, 112, 116, 130, 124, 116, 110, 109, 110, 105, 90, 89, 90, 101, 120, 122, 113, 116, 98, 95, 95, 84, 87, 91, 83, 101, 90, 79, 59, 55, 57, 65, 70, 82, 107, 104, 105, 113, 114, 110, 97, 84, 101, 115, 115, 104, 143, 139, 113, 101, 96, 117, 103, 106, 103, 99, 93, 111, 96, 94, 92, 130, 132, 77, 81, 96, 90, 85, 88, 102, 122, 103, 105, 106, 102, 97, 100, 96, 95, 93, 95, 98, 82, 103, 102, 107, 98, 98, 101, 102, 99, 104, 76, 98, 114, 109, 115, 100, 90, 81, 44, 73, 50, 100, 135, 120, 120, 115, 112, 114, 117, 125, 125, 123, 129, 136, 127, 120, 125, 128, 123, 137, 146, 134, 126, 127, 122, 141, 129, 131, 123, 121, 83, 91, 156, 150, 102, 104, 128, 139, 139, 135, 155, 145, 150, 145, 158, 154, 148, 132, 156, 166, 178, 161, 157, 151, 154, 162, 166, 163, 168, 167, 175, 164, 163, 165, 165, 137, 137, 133, 125, 145, 136, 138, 136, 132, 127, 138, 132, 138, 135, 128, 126, 120, 126, 129, 139, 125, 122, 127, 130, 130, 115, 118, 120, 126, 120, 120, 119, 116, 144, 160, 127, 117, 135, 116, 141, 123, 121, 136, 132, 128, 136, 133, 132, 132, 134, 127, 132, 134, 124, 123, 124, 128, 127, 116, 120, 114, 117, 118, 125, 123, 123, 120, 107, 115, 103, 99, 105, 104, 109, 110, 109, 108, 95, 106, 108, 99, 103, 102, 105, 112, 126, 120, 119, 113, 116, 118, 126, 141, 128, 120, 118, 111, 103, 103, 94, 95, 101, 100, 111, 120, 112, 97, 97, 100, 96, 93, 97, 99, 87, 92, 84, 76, 60, 58, 55, 64, 78, 92, 111, 101, 112, 111, 111, 111, 101, 96, 100, 116, 102, 82, 111, 119, 118, 102, 100, 116, 102, 106, 110, 106, 93, 112, 74, 62, 100, 128, 157, 159, 88, 92, 89, 82, 98, 94, 111, 101, 108, 101, 105, 77, 98, 93, 95, 94, 91, 95, 88, 105, 103, 107, 104, 98, 96, 105, 102, 104, 102, 105, 118, 107, 102, 103, 92, 85, 61, 69, 70, 81, 119, 123, 126, 113, 110, 109, 120, 123, 129, 128, 128, 131, 124, 132, 131, 126, 131, 148, 139, 128, 126, 126, 116, 136, 127, 118, 116, 121, 78, 69, 111, 132, 131, 125, 140, 136, 142, 137, 154, 151, 148, 146, 155, 151, 149, 137, 149, 168, 168, 156, 157, 159, 160, 165, 158, 153, 158, 168, 160, 169, 166, 166, 164, 135, 139, 132, 123, 127, 142, 125, 144, 139, 128, 136, 133, 127, 128, 133, 128, 111, 142, 140, 126, 137, 117, 119, 132, 126, 124, 127, 138, 127, 110, 130, 95, 105, 135, 154, 120, 124, 130, 132, 142, 127, 127, 134, 135, 131, 127, 129, 132, 128, 134, 124, 127, 131, 126, 127, 121, 133, 126, 123, 132, 131, 115, 123, 127, 129, 120, 119, 119, 110, 119, 114, 108, 107, 118, 120, 107, 118, 116, 119, 113, 104, 95, 104, 115, 116, 118, 111, 105, 100, 119, 119, 141, 135, 130, 123, 119, 106, 85, 93, 91, 97, 99, 98, 105, 109, 104, 92, 79, 82, 101, 99, 94, 92, 96, 92, 87, 71, 57, 57, 51, 58, 69, 81, 109, 104, 108, 109, 107, 113, 100, 104, 107, 115, 111, 97, 102, 89, 123, 113, 104, 117, 107, 108, 108, 109, 105, 91, 58, 68, 94, 138, 164, 185, 115, 92, 89, 89, 109, 110, 102, 107, 104, 105, 101, 112, 102, 101, 92, 106, 89, 84, 96, 102, 98, 108, 102, 101, 106, 104, 104, 103, 112, 110, 132, 119, 115, 109, 101, 109, 93, 86, 91, 88, 105, 115, 124, 115, 112, 101, 118, 123, 132, 127, 131, 130, 128, 127, 132, 130, 131, 133, 134, 138, 124, 125, 128, 129, 128, 124, 123, 107, 104, 89, 82, 96, 112, 134, 148, 144, 146, 146, 150, 149, 152, 153, 155, 148, 158, 150, 145, 144, 165, 156, 169, 158, 143, 159, 157, 155, 166, 173, 167, 169, 167, 169, 166, 136, 140, 134, 133, 116, 130, 125, 133, 127, 143, 127, 130, 130, 132, 129, 134, 105, 135, 130, 117, 147, 132, 137, 133, 122, 138, 132, 140, 120, 109, 143, 147, 115, 127, 127, 129, 131, 127, 131, 145, 139, 130, 134, 135, 124, 129, 142, 130, 128, 126, 121, 131, 118, 131, 142, 133, 127, 126, 126, 128, 121, 125, 128, 127, 121, 117, 120, 115, 106, 119, 113, 110, 111, 93, 105, 101, 108, 108, 119, 99, 106, 105, 106, 112, 117, 121, 108, 113, 116, 118, 125, 145, 131, 122, 119, 114, 108, 90, 87, 85, 91, 94, 97, 96, 90, 96, 91, 89, 85, 93, 101, 99, 97, 98, 91, 85, 63, 47, 41, 43, 45, 56, 77, 95, 99, 96, 105, 123, 110, 106, 119, 112, 114, 119, 105, 110, 94, 101, 130, 111, 108, 105, 105, 102, 107, 98, 82, 51, 67, 88, 133, 155, 156, 99, 122, 107, 109, 103, 103, 107, 110, 112, 112, 96, 105, 108, 96, 101, 104, 102, 96, 100, 104, 102, 105, 108, 97, 110, 106, 113, 105, 108, 119, 128, 128, 122, 112, 108, 114, 106, 102, 103, 96, 102, 115, 129, 114, 107, 115, 117, 124, 128, 121, 132, 129, 127, 124, 131, 119, 130, 126, 128, 112, 139, 122, 128, 123, 131, 129, 118, 115, 108, 93, 89, 104, 121, 132, 143, 151, 151, 152, 159, 152, 153, 147, 149, 151, 156, 154, 151, 151, 157, 157, 162, 162, 150, 161, 158, 149, 165, 168, 163, 163, 163, 161, 160, 137, 138, 119, 133, 124, 141, 131, 138, 135, 136, 128, 127, 123, 120, 137, 135, 133, 132, 125, 125, 130, 152, 131, 142, 133, 128, 136, 135, 131, 94, 131, 152, 126, 139, 136, 117, 135, 145, 138, 142, 131, 137, 141, 131, 124, 131, 124, 120, 136, 130, 124, 117, 91, 130, 140, 123, 134, 126, 124, 118, 130, 121, 131, 113, 119, 104, 115, 110, 115, 114, 107, 115, 115, 108, 105, 116, 114, 91, 107, 105, 113, 109, 111, 120, 118, 119, 102, 107, 116, 118, 137, 149, 138, 121, 129, 122, 107, 83, 81, 80, 89, 89, 93, 91, 91, 86, 96, 87, 88, 99, 92, 106, 108, 101, 98, 90, 62, 52, 31, 7, 24, 46, 71, 90, 96, 103, 106, 114, 111, 112, 104, 112, 114, 119, 114, 98, 104, 105, 113, 106, 106, 106, 85, 89, 99, 92, 78, 48, 69, 94, 120, 138, 142, 84, 98, 119, 115, 99, 110, 111, 104, 115, 112, 110, 112, 109, 93, 94, 105, 102, 102, 100, 118, 102, 108, 105, 113, 110, 106, 116, 110, 114, 116, 115, 130, 106, 120, 110, 124, 114, 110, 103, 112, 105, 114, 119, 112, 110, 115, 104, 121, 126, 117, 120, 125, 126, 124, 127, 121, 131, 130, 132, 121, 116, 132, 133, 125, 122, 123, 118, 113, 112, 102, 105, 109, 125, 140, 142, 152, 152, 149, 158, 155, 150, 152, 154, 158, 154, 156, 159, 154, 159, 160, 155, 159, 154, 164, 158, 158, 165, 164, 164, 163, 167, 167, 173, 136, 145, 132, 132, 141, 131, 133, 137, 147, 138, 137, 132, 136, 137, 132, 109, 128, 135, 144, 128, 131, 140, 141, 136, 130, 134, 131, 124, 143, 128, 139, 130, 118, 139, 104, 124, 122, 143, 139, 128, 136, 134, 127, 141, 138, 126, 128, 113, 126, 145, 127, 123, 102, 121, 140, 126, 120, 126, 126, 124, 130, 130, 123, 129, 126, 105, 125, 108, 119, 121, 118, 120, 120, 106, 110, 110, 104, 103, 113, 115, 106, 104, 116, 112, 113, 116, 97, 107, 119, 119, 147, 151, 141, 142, 137, 131, 103, 92, 86, 83, 87, 86, 89, 80, 89, 76, 91, 93, 95, 93, 99, 96, 94, 98, 93, 82, 64, 51, 21, 0, 12, 42, 71, 86, 94, 101, 113, 117, 114, 105, 113, 111, 111, 107, 115, 109, 106, 106, 111, 107, 101, 80, 76, 66, 82, 89, 86, 61, 57, 79, 107, 127, 120, 96, 85, 111, 106, 110, 119, 106, 82, 112, 113, 108, 105, 107, 108, 101, 106, 103, 110, 109, 103, 114, 115, 111, 112, 111, 116, 109, 109, 107, 116, 115, 123, 111, 123, 100, 125, 114, 117, 108, 117, 116, 108, 111, 118, 118, 115, 99, 117, 115, 112, 122, 124, 126, 115, 125, 138, 134, 130, 126, 126, 116, 136, 129, 125, 127, 121, 114, 115, 116, 112, 118, 115, 137, 146, 144, 150, 156, 149, 152, 153, 148, 153, 147, 151, 154, 155, 150, 154, 160, 156, 157, 159, 158, 159, 164, 161, 165, 162, 159, 163, 160, 161, 169, 141, 138, 129, 128, 129, 122, 126, 145, 145, 128, 136, 139, 138, 128, 134, 129, 133, 136, 133, 134, 135, 131, 139, 136, 142, 129, 126, 140, 137, 125, 139, 140, 130, 126, 130, 119, 115, 136, 132, 140, 129, 125, 132, 132, 141, 136, 132, 113, 130, 128, 118, 133, 117, 112, 125, 122, 119, 127, 128, 136, 134, 127, 131, 131, 130, 112, 125, 122, 116, 114, 106, 109, 113, 106, 102, 110, 111, 101, 98, 112, 110, 99, 108, 108, 111, 114, 111, 118, 119, 124, 146, 140, 146, 149, 132, 129, 100, 95, 97, 89, 90, 88, 80, 85, 83, 86, 93, 91, 93, 90, 90, 89, 83, 88, 95, 87, 60, 50, 32, 21, 29, 52, 78, 94, 97, 106, 93, 118, 115, 124, 113, 114, 116, 115, 114, 114, 110, 107, 110, 101, 97, 82, 56, 58, 83, 103, 91, 91, 71, 76, 92, 107, 92, 94, 106, 111, 98, 115, 120, 114, 106, 109, 113, 110, 116, 111, 111, 106, 106, 104, 104, 105, 108, 110, 105, 104, 109, 107, 109, 92, 103, 103, 110, 110, 115, 115, 117, 119, 119, 123, 124, 114, 122, 119, 111, 106, 122, 118, 115, 102, 106, 115, 117, 125, 117, 130, 100, 120, 141, 130, 123, 125, 122, 127, 129, 128, 127, 125, 127, 117, 116, 116, 136, 113, 114, 157, 156, 147, 143, 143, 150, 151, 152, 150, 151, 145, 145, 149, 140, 144, 152, 154, 156, 157, 158, 160, 161, 153, 161, 165, 167, 170, 164, 167, 164, 175, 127, 125, 118, 129, 129, 124, 129, 135, 134, 130, 138, 139, 142, 138, 139, 139, 141, 147, 123, 126, 136, 135, 140, 144, 128, 147, 143, 133, 127, 108, 133, 128, 139, 128, 143, 131, 131, 123, 126, 149, 131, 129, 130, 131, 127, 129, 140, 129, 125, 120, 118, 126, 133, 133, 122, 123, 135, 128, 128, 129, 131, 129, 134, 123, 123, 102, 118, 132, 114, 97, 120, 114, 101, 111, 105, 112, 98, 89, 98, 111, 108, 100, 112, 116, 114, 112, 111, 112, 111, 118, 151, 139, 143, 148, 138, 134, 113, 110, 102, 95, 88, 94, 87, 87, 83, 94, 98, 86, 93, 91, 90, 88, 91, 93, 94, 87, 70, 55, 35, 40, 51, 60, 84, 88, 95, 103, 107, 106, 102, 110, 116, 115, 112, 112, 116, 122, 110, 107, 99, 118, 122, 93, 82, 86, 95, 101, 105, 107, 100, 87, 93, 104, 101, 90, 101, 117, 108, 112, 113, 122, 107, 109, 112, 108, 110, 107, 103, 110, 110, 109, 107, 99, 106, 110, 109, 106, 109, 105, 109, 106, 105, 112, 108, 112, 120, 118, 128, 124, 124, 118, 107, 116, 121, 137, 112, 100, 112, 105, 101, 97, 98, 101, 113, 129, 127, 128, 118, 124, 129, 118, 124, 124, 126, 135, 118, 121, 129, 124, 122, 120, 118, 111, 130, 108, 123, 142, 152, 149, 155, 144, 155, 155, 152, 153, 152, 152, 144, 153, 148, 155, 155, 160, 160, 162, 163, 147, 157, 157, 157, 167, 165, 162, 163, 151, 180, 162, 132, 121, 119, 119, 138, 133, 137, 137, 128, 142, 139, 144, 138, 135, 136, 132, 140, 137, 136, 139, 134, 134, 138, 137, 122, 143, 125, 137, 164, 125, 143, 135, 123, 140, 124, 139, 139, 129, 128, 137, 125, 132, 124, 141, 128, 138, 133, 125, 102, 118, 124, 119, 141, 136, 129, 132, 129, 130, 129, 128, 142, 126, 120, 127, 129, 122, 131, 126, 110, 96, 94, 95, 114, 117, 112, 108, 95, 90, 113, 100, 124, 107, 120, 121, 116, 108, 113, 115, 116, 122, 143, 139, 146, 152, 143, 141, 122, 109, 103, 98, 92, 94, 91, 94, 86, 89, 92, 89, 89, 98, 98, 92, 101, 89, 93, 86, 68, 60, 36, 56, 73, 71, 76, 82, 93, 98, 115, 103, 107, 100, 113, 114, 109, 112, 107, 111, 110, 90, 100, 120, 139, 118, 102, 104, 105, 102, 116, 108, 108, 103, 105, 104, 109, 100, 106, 116, 115, 113, 112, 116, 100, 113, 111, 113, 108, 108, 111, 112, 109, 109, 113, 92, 106, 98, 105, 116, 107, 105, 111, 109, 107, 106, 106, 115, 122, 115, 127, 122, 123, 90, 113, 103, 123, 145, 134, 107, 107, 106, 103, 86, 74, 85, 113, 119, 122, 125, 129, 128, 130, 120, 124, 125, 124, 126, 126, 122, 133, 130, 119, 117, 124, 122, 124, 130, 130, 139, 139, 149, 146, 154, 147, 148, 154, 153, 151, 153, 147, 151, 158, 158, 153, 153, 156, 162, 160, 156, 153, 166, 151, 162, 160, 166, 165, 162, 163, 168, 131, 133, 130, 134, 128, 126, 138, 136, 136, 137, 142, 146, 138, 136, 141, 141, 134, 133, 141, 140, 137, 131, 138, 139, 132, 133, 93, 135, 174, 160, 138, 132, 125, 136, 130, 137, 134, 126, 132, 135, 126, 125, 130, 133, 131, 137, 134, 129, 121, 123, 144, 125, 129, 127, 127, 131, 127, 131, 131, 129, 132, 122, 126, 127, 126, 129, 127, 109, 128, 123, 104, 112, 107, 120, 119, 110, 103, 107, 113, 109, 107, 109, 123, 97, 110, 111, 109, 115, 105, 110, 127, 129, 146, 156, 151, 140, 131, 120, 109, 107, 104, 99, 98, 98, 99, 95, 86, 82, 78, 81, 92, 94, 99, 93, 89, 80, 79, 50, 41, 66, 70, 76, 66, 63, 77, 96, 113, 104, 103, 98, 103, 107, 100, 108, 114, 94, 116, 85, 104, 116, 127, 119, 112, 95, 107, 96, 102, 100, 105, 108, 108, 102, 115, 110, 111, 107, 113, 117, 109, 119, 107, 122, 109, 107, 113, 115, 113, 112, 115, 103, 111, 108, 104, 90, 105, 121, 102, 120, 114, 112, 111, 118, 104, 121, 116, 120, 122, 124, 116, 105, 113, 103, 112, 138, 130, 115, 102, 104, 100, 75, 41, 74, 104, 112, 118, 120, 119, 123, 133, 126, 131, 121, 125, 126, 124, 130, 115, 131, 133, 125, 126, 127, 126, 134, 146, 141, 146, 145, 135, 154, 149, 146, 153, 154, 150, 150, 148, 159, 155, 153, 143, 155, 156, 155, 154, 167, 159, 159, 155, 170, 148, 160, 164, 170, 164, 163, 134, 130, 128, 134, 130, 134, 141, 134, 137, 132, 138, 140, 127, 147, 133, 143, 138, 142, 133, 145, 118, 137, 162, 139, 130, 135, 114, 119, 145, 142, 142, 136, 130, 136, 137, 133, 147, 125, 137, 137, 125, 131, 134, 132, 129, 130, 131, 118, 135, 133, 135, 134, 126, 122, 137, 126, 133, 129, 130, 124, 131, 115, 118, 136, 123, 130, 122, 93, 131, 146, 131, 111, 98, 101, 114, 106, 112, 111, 107, 102, 109, 106, 118, 113, 111, 113, 100, 116, 109, 123, 143, 134, 137, 159, 157, 147, 138, 124, 118, 109, 102, 96, 104, 98, 101, 94, 82, 85, 72, 80, 90, 86, 80, 76, 75, 75, 72, 62, 50, 56, 65, 75, 65, 52, 73, 94, 101, 102, 99, 96, 79, 95, 108, 110, 109, 117, 114, 102, 103, 112, 124, 104, 96, 103, 101, 104, 105, 99, 103, 112, 107, 107, 113, 111, 102, 108, 109, 120, 117, 121, 115, 122, 109, 103, 99, 114, 112, 108, 121, 114, 110, 109, 104, 83, 110, 118, 105, 112, 115, 121, 124, 131, 107, 130, 112, 117, 129, 123, 116, 116, 113, 111, 113, 118, 113, 120, 102, 108, 107, 95, 66, 75, 95, 116, 112, 122, 119, 124, 126, 133, 136, 125, 112, 114, 125, 123, 116, 123, 134, 120, 135, 126, 130, 140, 139, 138, 127, 161, 148, 146, 152, 148, 139, 151, 158, 156, 149, 154, 139, 172, 167, 154, 157, 148, 162, 156, 165, 160, 163, 161, 163, 158, 164, 165, 162, 176, 141, 132, 128, 141, 136, 131, 136, 139, 136, 132, 138, 132, 138, 139, 138, 141, 138, 137, 129, 144, 121, 131, 150, 141, 144, 138, 125, 136, 136, 139, 142, 140, 142, 131, 137, 136, 145, 135, 130, 128, 132, 135, 130, 140, 133, 123, 138, 129, 132, 138, 131, 135, 133, 132, 136, 133, 125, 121, 130, 127, 132, 120, 123, 133, 132, 128, 117, 91, 102, 135, 148, 116, 100, 94, 110, 102, 108, 108, 100, 109, 112, 111, 105, 121, 115, 111, 107, 111, 111, 117, 139, 140, 137, 151, 163, 160, 142, 127, 119, 104, 95, 90, 118, 108, 108, 90, 85, 94, 88, 83, 86, 78, 73, 69, 79, 73, 71, 62, 62, 55, 52, 67, 66, 48, 67, 82, 94, 107, 104, 96, 91, 94, 105, 109, 106, 113, 107, 110, 112, 114, 119, 113, 98, 105, 104, 107, 113, 111, 100, 110, 113, 114, 114, 118, 113, 101, 114, 104, 108, 115, 105, 111, 116, 114, 115, 108, 108, 109, 109, 113, 110, 114, 108, 107, 93, 105, 109, 115, 112, 119, 120, 125, 120, 117, 120, 114, 127, 121, 136, 103, 115, 114, 117, 112, 113, 111, 116, 118, 112, 116, 107, 98, 114, 114, 109, 128, 123, 126, 128, 131, 130, 127, 125, 134, 126, 128, 131, 134, 129, 122, 124, 123, 130, 139, 147, 137, 133, 162, 145, 141, 146, 149, 147, 151, 159, 153, 148, 145, 120, 164, 169, 160, 152, 162, 150, 154, 157, 167, 161, 163, 165, 163, 165, 168, 169, 167, 132, 145, 134, 130, 142, 131, 146, 138, 139, 132, 136, 137, 141, 140, 137, 129, 131, 144, 129, 137, 137, 131, 133, 137, 132, 143, 133, 139, 147, 131, 138, 137, 144, 134, 139, 137, 147, 136, 133, 143, 132, 141, 126, 134, 127, 134, 137, 131, 125, 137, 140, 137, 135, 136, 137, 135, 132, 125, 125, 125, 115, 127, 130, 129, 128, 119, 140, 101, 103, 119, 102, 104, 107, 109, 112, 111, 99, 107, 117, 112, 116, 113, 111, 111, 109, 117, 115, 111, 105, 116, 143, 147, 144, 151, 157, 165, 140, 124, 124, 114, 100, 94, 99, 104, 107, 106, 104, 107, 98, 90, 86, 72, 61, 63, 68, 72, 64, 52, 49, 61, 69, 72, 63, 49, 64, 75, 77, 93, 106, 100, 96, 101, 101, 100, 105, 112, 112, 109, 108, 115, 113, 114, 108, 105, 105, 108, 118, 117, 115, 116, 96, 95, 117, 153, 160, 106, 116, 99, 101, 106, 98, 113, 107, 102, 109, 106, 114, 114, 111, 109, 112, 114, 108, 112, 93, 107, 114, 114, 112, 118, 121, 120, 123, 110, 128, 117, 129, 129, 132, 126, 121, 118, 102, 103, 114, 110, 112, 119, 122, 124, 116, 118, 118, 123, 128, 126, 117, 132, 135, 130, 134, 134, 130, 135, 124, 132, 136, 138, 127, 119, 133, 133, 136, 135, 139, 146, 141, 151, 142, 143, 156, 157, 149, 149, 155, 158, 155, 157, 157, 153, 157, 157, 161, 155, 161, 165, 164, 163, 168, 163, 170, 160, 168, 167, 161, 167, 133, 140, 132, 133, 143, 134, 132, 136, 141, 128, 142, 139, 134, 126, 130, 138, 139, 137, 124, 143, 136, 136, 138, 134, 130, 139, 135, 137, 139, 142, 135, 148, 143, 131, 130, 143, 137, 143, 132, 140, 139, 130, 130, 128, 126, 151, 135, 129, 137, 134, 133, 137, 127, 138, 131, 135, 126, 117, 133, 133, 135, 127, 124, 125, 127, 126, 126, 115, 120, 119, 108, 113, 118, 114, 106, 102, 103, 103, 113, 107, 112, 110, 115, 107, 107, 111, 116, 113, 112, 127, 146, 158, 145, 155, 160, 173, 148, 116, 128, 114, 109, 103, 109, 116, 114, 102, 108, 110, 108, 94, 82, 74, 52, 54, 61, 65, 66, 68, 68, 66, 81, 81, 66, 53, 67, 74, 69, 73, 92, 102, 98, 103, 108, 98, 103, 113, 116, 114, 111, 114, 120, 115, 107, 108, 110, 110, 110, 113, 115, 118, 71, 71, 106, 152, 187, 119, 117, 111, 108, 111, 107, 107, 108, 104, 103, 112, 108, 110, 111, 113, 112, 108, 104, 102, 99, 111, 114, 117, 117, 109, 115, 122, 125, 118, 122, 129, 140, 137, 136, 124, 116, 114, 104, 106, 113, 115, 114, 111, 122, 120, 121, 124, 124, 125, 133, 124, 128, 132, 136, 148, 138, 135, 129, 126, 126, 133, 137, 137, 129, 127, 130, 133, 140, 135, 140, 149, 142, 152, 144, 145, 153, 154, 148, 146, 152, 157, 155, 156, 157, 158, 164, 153, 154, 160, 159, 168, 162, 156, 156, 163, 167, 165, 158, 170, 170, 169, 151, 141, 126, 143, 139, 137, 140, 130, 144, 132, 136, 138, 134, 138, 134, 139, 137, 137, 143, 146, 139, 131, 131, 152, 142, 133, 136, 142, 134, 122, 146, 156, 136, 128, 144, 138, 109, 142, 143, 144, 142, 128, 127, 121, 126, 144, 134, 122, 110, 140, 131, 123, 120, 163, 145, 126, 112, 126, 137, 131, 135, 134, 126, 126, 127, 116, 119, 121, 118, 115, 123, 109, 109, 114, 112, 104, 104, 114, 109, 95, 112, 108, 110, 109, 110, 109, 109, 96, 89, 128, 141, 153, 148, 151, 158, 153, 147, 131, 123, 116, 113, 112, 114, 112, 98, 101, 110, 110, 104, 89, 78, 69, 63, 63, 65, 58, 56, 70, 68, 72, 80, 83, 65, 52, 53, 58, 62, 68, 77, 92, 97, 95, 106, 102, 104, 106, 111, 118, 112, 114, 113, 117, 114, 112, 97, 109, 115, 111, 108, 125, 67, 64, 107, 137, 157, 113, 113, 112, 110, 119, 113, 98, 103, 105, 109, 112, 113, 112, 110, 113, 115, 109, 104, 106, 102, 110, 106, 108, 123, 114, 114, 123, 123, 121, 131, 141, 148, 138, 125, 113, 109, 108, 102, 105, 105, 109, 110, 110, 123, 114, 130, 112, 123, 126, 136, 135, 129, 127, 138, 139, 131, 125, 134, 126, 132, 135, 132, 133, 133, 132, 137, 130, 135, 145, 136, 148, 150, 147, 144, 143, 146, 147, 157, 155, 154, 154, 150, 155, 155, 162, 148, 164, 162, 155, 158, 163, 157, 156, 169, 158, 154, 170, 161, 167, 174, 151, 142, 133, 126, 116, 136, 131, 137, 132, 138, 141, 140, 134, 143, 131, 134, 132, 141, 147, 137, 138, 139, 124, 138, 143, 138, 140, 138, 146, 140, 118, 141, 165, 138, 140, 143, 136, 120, 132, 140, 146, 141, 135, 138, 134, 128, 121, 129, 134, 114, 129, 138, 132, 111, 146, 132, 110, 122, 116, 126, 125, 124, 122, 129, 129, 121, 116, 125, 123, 121, 127, 119, 111, 114, 112, 105, 106, 105, 113, 107, 102, 100, 114, 113, 108, 106, 110, 117, 108, 100, 136, 146, 156, 149, 153, 160, 148, 149, 152, 131, 122, 113, 118, 106, 108, 105, 108, 110, 109, 90, 88, 84, 55, 61, 49, 50, 51, 49, 61, 70, 80, 87, 87, 71, 60, 65, 55, 70, 68, 71, 79, 88, 92, 88, 103, 110, 114, 111, 115, 115, 113, 111, 111, 116, 123, 110, 109, 111, 119, 117, 136, 85, 64, 94, 129, 118, 106, 125, 104, 87, 120, 141, 107, 105, 107, 106, 113, 113, 116, 113, 118, 112, 109, 108, 115, 115, 103, 104, 113, 113, 116, 119, 127, 123, 131, 132, 141, 144, 141, 128, 121, 108, 109, 105, 114, 112, 114, 117, 114, 116, 108, 125, 117, 111, 133, 142, 141, 132, 132, 138, 136, 122, 126, 123, 129, 129, 125, 135, 133, 138, 131, 124, 132, 135, 141, 146, 140, 147, 154, 153, 146, 153, 158, 156, 145, 149, 156, 156, 153, 155, 150, 139, 168, 193, 150, 161, 150, 161, 162, 161, 171, 159, 174, 168, 167, 165, 168, 139, 135, 147, 109, 118, 117, 129, 129, 141, 133, 139, 124, 137, 145, 137, 133, 140, 133, 138, 137, 135, 131, 132, 140, 142, 144, 141, 140, 139, 131, 131, 144, 141, 131, 145, 137, 127, 125, 133, 130, 140, 130, 138, 124, 131, 137, 126, 127, 133, 130, 131, 133, 121, 134, 129, 132, 139, 131, 120, 120, 127, 132, 136, 123, 136, 116, 122, 123, 119, 116, 109, 116, 117, 116, 115, 104, 113, 105, 113, 113, 114, 107, 120, 120, 101, 116, 113, 102, 120, 145, 146, 149, 146, 142, 156, 152, 147, 151, 141, 128, 124, 128, 117, 115, 118, 114, 114, 109, 89, 83, 101, 69, 62, 54, 42, 40, 45, 51, 70, 82, 85, 75, 63, 62, 66, 61, 64, 70, 65, 70, 81, 93, 90, 91, 99, 107, 112, 110, 116, 111, 112, 112, 98, 125, 100, 111, 106, 114, 112, 126, 97, 81, 92, 103, 99, 106, 119, 106, 85, 117, 131, 111, 93, 104, 130, 116, 113, 115, 112, 115, 116, 115, 115, 111, 104, 112, 112, 116, 119, 117, 121, 124, 124, 128, 128, 140, 144, 141, 131, 123, 111, 108, 107, 85, 110, 120, 116, 117, 119, 113, 127, 119, 123, 126, 133, 146, 139, 129, 139, 140, 118, 120, 125, 135, 121, 128, 131, 131, 129, 127, 125, 135, 139, 145, 140, 146, 143, 150, 153, 145, 149, 155, 151, 147, 152, 158, 155, 154, 151, 151, 131, 163, 178, 154, 170, 161, 162, 159, 156, 167, 173, 167, 165, 169, 171, 164, 134, 136, 138, 127, 131, 123, 139, 128, 143, 134, 141, 118, 111, 142, 134, 137, 144, 139, 142, 131, 136, 137, 129, 137, 135, 142, 136, 146, 147, 138, 145, 145, 144, 134, 138, 142, 138, 138, 140, 136, 135, 136, 146, 132, 136, 134, 130, 125, 138, 132, 130, 132, 141, 137, 136, 135, 137, 129, 129, 128, 126, 133, 120, 118, 129, 121, 121, 124, 116, 114, 116, 109, 94, 106, 111, 119, 114, 105, 108, 107, 109, 122, 113, 117, 114, 105, 117, 116, 113, 139, 143, 137, 141, 143, 146, 149, 149, 145, 139, 127, 123, 113, 127, 125, 122, 107, 106, 101, 99, 83, 73, 54, 63, 55, 46, 41, 52, 59, 61, 71, 88, 75, 58, 64, 61, 61, 61, 65, 69, 75, 75, 78, 83, 91, 90, 96, 103, 114, 115, 112, 112, 113, 110, 108, 96, 107, 106, 107, 107, 111, 95, 96, 93, 90, 101, 103, 113, 113, 94, 104, 102, 91, 72, 101, 138, 133, 110, 117, 118, 120, 118, 119, 114, 113, 112, 111, 115, 114, 119, 120, 117, 111, 105, 121, 126, 142, 139, 140, 135, 124, 113, 107, 101, 89, 93, 115, 120, 116, 126, 122, 128, 123, 130, 137, 135, 139, 129, 130, 136, 129, 126, 133, 129, 122, 126, 132, 127, 129, 123, 125, 128, 138, 141, 148, 144, 147, 146, 149, 153, 140, 149, 155, 148, 155, 144, 149, 148, 154, 153, 153, 147, 158, 156, 148, 159, 170, 146, 166, 149, 157, 182, 175, 160, 162, 155, 166, 137, 133, 134, 135, 139, 118, 150, 142, 126, 140, 139, 125, 121, 135, 132, 138, 139, 148, 138, 131, 137, 129, 140, 138, 140, 134, 137, 133, 149, 133, 145, 131, 161, 143, 141, 146, 137, 147, 143, 137, 130, 139, 140, 133, 128, 133, 128, 129, 128, 139, 134, 127, 136, 136, 136, 137, 135, 131, 135, 124, 133, 123, 126, 127, 120, 117, 116, 106, 118, 122, 123, 115, 106, 112, 112, 113, 103, 118, 119, 111, 112, 115, 117, 113, 109, 115, 113, 132, 128, 139, 141, 139, 141, 140, 141, 132, 153, 143, 138, 127, 124, 90, 121, 125, 130, 112, 103, 108, 101, 85, 63, 57, 60, 61, 68, 58, 54, 61, 64, 78, 89, 81, 63, 55, 67, 70, 63, 58, 61, 69, 69, 65, 65, 81, 88, 106, 97, 100, 110, 106, 110, 108, 114, 100, 100, 102, 117, 106, 102, 108, 90, 93, 114, 106, 105, 94, 100, 123, 104, 101, 108, 100, 78, 91, 123, 114, 108, 115, 115, 122, 115, 122, 111, 108, 112, 98, 117, 111, 116, 118, 120, 89, 93, 121, 132, 138, 145, 143, 145, 129, 120, 107, 102, 98, 89, 108, 113, 110, 126, 120, 118, 117, 126, 134, 135, 128, 122, 133, 133, 124, 127, 137, 135, 132, 131, 126, 126, 128, 125, 126, 139, 137, 142, 144, 140, 154, 149, 151, 150, 153, 147, 152, 158, 156, 142, 145, 147, 152, 161, 161, 154, 162, 165, 155, 144, 179, 155, 167, 155, 153, 174, 155, 159, 169, 166, 171, 136, 128, 138, 140, 143, 136, 127, 107, 116, 140, 174, 169, 124, 129, 136, 129, 142, 140, 128, 131, 132, 135, 145, 142, 134, 134, 143, 143, 142, 138, 146, 132, 152, 139, 145, 138, 120, 149, 151, 144, 134, 140, 132, 134, 135, 135, 135, 131, 136, 129, 138, 133, 127, 130, 126, 137, 138, 130, 124, 128, 135, 136, 120, 119, 105, 120, 145, 106, 109, 112, 112, 120, 110, 91, 95, 120, 115, 115, 117, 114, 111, 114, 110, 120, 123, 128, 122, 137, 139, 139, 135, 141, 135, 136, 150, 134, 141, 155, 145, 126, 130, 128, 113, 118, 132, 113, 103, 108, 90, 85, 65, 61, 64, 64, 56, 61, 58, 67, 76, 71, 69, 84, 69, 58, 67, 71, 50, 48, 62, 69, 69, 59, 58, 68, 97, 105, 109, 110, 113, 114, 109, 105, 105, 106, 107, 104, 101, 106, 89, 102, 100, 101, 111, 102, 114, 97, 93, 127, 106, 104, 112, 109, 96, 106, 117, 105, 107, 115, 117, 117, 115, 122, 115, 116, 120, 115, 114, 119, 114, 116, 108, 108, 116, 128, 127, 130, 143, 146, 148, 130, 127, 100, 105, 95, 107, 120, 123, 119, 118, 126, 126, 121, 134, 127, 121, 135, 127, 128, 130, 121, 130, 139, 138, 128, 130, 126, 132, 123, 133, 132, 136, 135, 137, 148, 145, 145, 145, 153, 154, 149, 148, 146, 152, 150, 152, 149, 153, 155, 158, 159, 158, 158, 165, 164, 147, 159, 151, 165, 168, 162, 170, 157, 156, 163, 167, 172, 132, 135, 138, 142, 143, 149, 113, 82, 110, 138, 179, 208, 137, 130, 138, 124, 143, 146, 119, 134, 142, 137, 147, 140, 148, 121, 123, 175, 137, 138, 143, 138, 144, 144, 136, 137, 129, 145, 128, 146, 134, 139, 133, 132, 131, 123, 132, 134, 125, 128, 130, 134, 132, 130, 129, 122, 136, 123, 133, 126, 130, 126, 126, 94, 91, 157, 150, 118, 111, 114, 122, 122, 121, 113, 103, 118, 128, 118, 112, 116, 114, 115, 115, 102, 114, 138, 135, 137, 150, 141, 134, 132, 139, 137, 141, 135, 132, 139, 144, 136, 128, 129, 119, 113, 110, 110, 109, 115, 101, 71, 65, 58, 51, 52, 56, 66, 65, 62, 68, 69, 87, 88, 78, 73, 59, 64, 60, 48, 61, 66, 65, 66, 75, 74, 84, 109, 110, 113, 93, 135, 119, 109, 109, 111, 106, 103, 105, 100, 100, 103, 99, 97, 108, 105, 108, 100, 98, 111, 101, 105, 111, 111, 99, 107, 116, 114, 107, 101, 112, 116, 117, 113, 122, 116, 116, 112, 112, 125, 119, 118, 119, 124, 120, 133, 126, 131, 147, 145, 150, 136, 129, 106, 106, 95, 118, 123, 125, 115, 112, 110, 118, 124, 124, 135, 131, 128, 127, 131, 136, 119, 131, 136, 130, 121, 126, 133, 125, 134, 125, 136, 155, 136, 135, 138, 146, 136, 142, 148, 155, 143, 154, 148, 167, 142, 145, 146, 153, 156, 163, 161, 158, 151, 162, 160, 159, 158, 157, 157, 172, 162, 166, 155, 171, 167, 161, 169, 134, 138, 137, 138, 142, 147, 93, 76, 105, 134, 158, 202, 146, 129, 137, 136, 140, 137, 131, 139, 141, 140, 135, 143, 143, 139, 114, 150, 132, 131, 141, 136, 148, 137, 128, 151, 135, 138, 141, 141, 141, 134, 134, 130, 127, 127, 133, 116, 125, 123, 129, 142, 134, 132, 131, 137, 135, 128, 117, 125, 128, 119, 126, 85, 73, 166, 140, 114, 121, 123, 116, 117, 118, 104, 108, 108, 116, 112, 115, 93, 119, 123, 114, 111, 109, 125, 136, 137, 150, 145, 136, 141, 138, 134, 137, 142, 131, 129, 146, 133, 122, 119, 124, 117, 100, 95, 111, 111, 105, 89, 67, 59, 59, 52, 55, 63, 65, 71, 72, 72, 103, 101, 81, 82, 70, 57, 69, 55, 59, 63, 76, 74, 66, 76, 81, 103, 112, 106, 67, 126, 141, 122, 106, 105, 102, 109, 103, 98, 107, 109, 93, 102, 102, 90, 102, 100, 103, 111, 104, 104, 102, 106, 111, 113, 104, 108, 110, 99, 110, 112, 119, 114, 112, 118, 123, 119, 116, 118, 117, 120, 123, 123, 124, 126, 123, 130, 143, 141, 139, 131, 126, 124, 119, 118, 128, 123, 115, 116, 113, 101, 119, 127, 120, 133, 132, 124, 120, 134, 127, 113, 117, 131, 127, 126, 125, 127, 126, 136, 111, 132, 157, 138, 142, 136, 150, 139, 140, 145, 153, 147, 152, 138, 157, 140, 134, 152, 150, 164, 154, 158, 153, 166, 156, 162, 159, 156, 168, 167, 163, 164, 161, 165, 168, 161, 158, 165, 136, 136, 134, 134, 140, 142, 111, 77, 85, 125, 157, 181, 129, 126, 128, 142, 140, 139, 136, 143, 116, 136, 152, 121, 133, 151, 136, 142, 141, 141, 143, 134, 139, 140, 138, 141, 129, 144, 144, 141, 134, 134, 130, 133, 130, 131, 130, 127, 124, 132, 129, 134, 134, 129, 132, 133, 132, 122, 129, 124, 119, 118, 121, 124, 100, 122, 116, 105, 143, 123, 113, 124, 116, 111, 113, 111, 123, 116, 120, 120, 121, 119, 116, 119, 126, 137, 136, 141, 148, 140, 134, 140, 137, 138, 131, 128, 129, 130, 138, 134, 126, 118, 125, 123, 107, 108, 111, 115, 109, 87, 61, 59, 64, 59, 56, 59, 68, 66, 66, 80, 99, 108, 95, 87, 81, 60, 58, 55, 48, 65, 71, 74, 68, 70, 84, 102, 116, 112, 94, 97, 117, 110, 111, 108, 103, 96, 97, 102, 107, 109, 101, 102, 100, 98, 99, 91, 113, 110, 111, 99, 98, 109, 119, 118, 115, 117, 111, 116, 112, 109, 123, 121, 112, 114, 125, 118, 121, 117, 121, 118, 127, 128, 133, 120, 126, 130, 129, 139, 144, 135, 121, 130, 138, 136, 130, 124, 115, 114, 104, 109, 118, 124, 123, 126, 121, 104, 121, 128, 124, 117, 122, 124, 124, 131, 127, 128, 127, 126, 130, 134, 134, 129, 139, 140, 151, 133, 142, 148, 159, 142, 159, 143, 148, 152, 149, 153, 156, 150, 161, 164, 159, 165, 161, 162, 162, 152, 171, 157, 163, 167, 165, 160, 167, 168, 168, 161, 147, 137, 135, 137, 148, 145, 106, 106, 118, 104, 141, 139, 130, 129, 137, 140, 138, 146, 141, 134, 122, 128, 149, 137, 141, 140, 134, 140, 143, 139, 132, 130, 135, 145, 138, 143, 139, 141, 143, 130, 138, 138, 133, 133, 131, 118, 125, 128, 125, 122, 128, 130, 134, 123, 133, 132, 117, 129, 130, 121, 127, 126, 123, 125, 125, 126, 124, 92, 136, 113, 102, 121, 111, 106, 117, 104, 129, 115, 116, 112, 116, 115, 101, 125, 124, 138, 130, 133, 145, 129, 112, 132, 142, 139, 136, 132, 126, 122, 125, 132, 127, 114, 121, 112, 113, 103, 112, 106, 101, 83, 65, 55, 67, 63, 53, 66, 76, 68, 61, 82, 93, 101, 102, 97, 85, 72, 54, 58, 60, 56, 59, 68, 63, 75, 86, 103, 110, 110, 110, 115, 111, 95, 99, 103, 104, 99, 99, 97, 103, 108, 97, 103, 99, 97, 106, 106, 114, 109, 108, 104, 111, 104, 111, 114, 109, 114, 112, 114, 107, 103, 122, 105, 125, 110, 115, 113, 112, 112, 116, 118, 135, 136, 129, 119, 124, 116, 126, 132, 136, 133, 119, 130, 142, 131, 128, 121, 108, 106, 106, 112, 114, 122, 124, 123, 118, 92, 110, 125, 123, 119, 121, 123, 120, 136, 126, 130, 132, 115, 142, 135, 145, 136, 145, 137, 146, 149, 144, 150, 150, 139, 151, 152, 168, 159, 157, 153, 151, 147, 149, 154, 156, 154, 158, 161, 158, 151, 161, 154, 162, 158, 162, 156, 164, 163, 161, 167, 138, 143, 136, 143, 145, 129, 77, 149, 184, 123, 128, 129, 127, 139, 146, 137, 127, 162, 139, 134, 138, 137, 137, 140, 135, 142, 141, 133, 143, 134, 133, 127, 123, 142, 138, 137, 140, 143, 141, 133, 132, 127, 130, 139, 137, 129, 139, 127, 134, 128, 126, 131, 102, 129, 121, 128, 126, 122, 131, 134, 116, 130, 124, 121, 119, 131, 119, 117, 122, 119, 115, 121, 118, 114, 125, 118, 122, 113, 111, 113, 109, 108, 119, 115, 135, 135, 123, 139, 137, 117, 111, 134, 150, 145, 143, 140, 133, 120, 122, 129, 127, 120, 118, 115, 106, 108, 112, 114, 95, 73, 67, 70, 63, 61, 62, 64, 69, 70, 70, 94, 90, 90, 86, 87, 86, 75, 65, 66, 69, 59, 40, 57, 59, 73, 91, 99, 104, 105, 102, 114, 104, 102, 96, 108, 106, 104, 103, 105, 103, 103, 103, 106, 91, 96, 98, 106, 109, 108, 102, 102, 108, 102, 94, 112, 116, 114, 116, 110, 104, 110, 118, 103, 111, 108, 111, 97, 112, 117, 119, 120, 131, 135, 123, 120, 126, 122, 136, 123, 123, 123, 138, 146, 140, 139, 130, 123, 111, 102, 107, 112, 118, 124, 130, 124, 123, 124, 118, 122, 126, 125, 121, 120, 119, 131, 123, 115, 122, 125, 139, 132, 136, 150, 136, 141, 137, 150, 149, 147, 145, 145, 146, 149, 155, 154, 149, 156, 154, 157, 154, 156, 154, 145, 157, 157, 157, 157, 159, 148, 158, 162, 164, 160, 161, 164, 164, 169, 134, 142, 141, 137, 148, 123, 59, 140, 171, 114, 132, 131, 118, 129, 135, 134, 131, 141, 141, 139, 137, 132, 140, 138, 146, 138, 145, 139, 132, 137, 137, 139, 130, 138, 136, 136, 139, 141, 145, 138, 130, 132, 135, 140, 135, 130, 138, 122, 133, 135, 125, 132, 128, 122, 126, 122, 120, 126, 122, 120, 121, 131, 126, 127, 132, 122, 120, 117, 117, 120, 116, 117, 107, 116, 114, 126, 114, 118, 119, 115, 116, 111, 110, 129, 137, 129, 134, 145, 138, 137, 127, 141, 147, 141, 139, 141, 140, 124, 133, 133, 115, 115, 117, 113, 111, 116, 120, 117, 85, 73, 67, 74, 65, 62, 62, 76, 83, 84, 76, 78, 86, 84, 88, 86, 84, 75, 68, 63, 64, 52, 34, 49, 64, 78, 89, 101, 100, 107, 100, 106, 100, 97, 98, 99, 100, 96, 97, 97, 105, 107, 103, 101, 105, 101, 101, 108, 109, 107, 111, 108, 100, 103, 105, 102, 118, 104, 108, 108, 106, 117, 108, 108, 115, 107, 114, 99, 117, 119, 114, 125, 126, 125, 119, 105, 132, 138, 122, 127, 128, 130, 131, 147, 143, 138, 139, 129, 115, 111, 109, 113, 119, 114, 128, 122, 123, 134, 122, 114, 124, 117, 125, 116, 125, 126, 128, 122, 120, 131, 139, 137, 140, 145, 141, 142, 136, 146, 146, 154, 150, 149, 152, 156, 151, 153, 158, 148, 145, 151, 149, 163, 152, 150, 153, 154, 159, 162, 154, 153, 155, 161, 156, 155, 163, 159, 164, 169, 141, 144, 145, 137, 144, 138, 115, 128, 132, 124, 141, 121, 125, 116, 134, 142, 132, 135, 139, 134, 141, 139, 141, 140, 139, 130, 128, 138, 131, 128, 144, 139, 138, 133, 117, 139, 138, 140, 139, 132, 129, 132, 135, 138, 135, 134, 128, 121, 126, 122, 121, 123, 118, 121, 122, 125, 128, 124, 119, 132, 129, 118, 123, 100, 143, 120, 119, 120, 117, 114, 124, 118, 118, 123, 112, 124, 122, 115, 112, 118, 120, 112, 114, 122, 132, 137, 140, 155, 139, 137, 127, 147, 152, 149, 142, 147, 132, 132, 139, 131, 120, 111, 113, 118, 121, 121, 120, 115, 102, 77, 71, 77, 71, 63, 58, 61, 58, 79, 89, 75, 91, 90, 79, 82, 83, 77, 77, 61, 63, 48, 33, 40, 59, 70, 88, 99, 94, 104, 102, 98, 97, 105, 103, 104, 95, 100, 100, 101, 104, 104, 94, 111, 97, 99, 98, 105, 103, 108, 98, 109, 102, 98, 103, 87, 109, 106, 103, 101, 116, 106, 101, 94, 104, 109, 112, 121, 120, 109, 117, 135, 133, 129, 121, 120, 125, 134, 125, 120, 120, 122, 125, 143, 138, 141, 144, 135, 130, 122, 117, 108, 110, 116, 117, 121, 124, 128, 118, 118, 121, 127, 124, 122, 111, 123, 123, 119, 113, 128, 137, 137, 138, 138, 139, 147, 139, 141, 149, 153, 151, 145, 154, 148, 154, 152, 153, 149, 160, 155, 153, 159, 160, 147, 160, 158, 151, 157, 163, 151, 157, 158, 144, 158, 162, 157, 161, 168, 134, 155, 138, 134, 140, 136, 143, 135, 136, 134, 136, 121, 133, 135, 132, 139, 138, 137, 142, 135, 136, 134, 138, 146, 134, 134, 136, 124, 163, 124, 129, 136, 135, 142, 129, 137, 148, 133, 136, 140, 130, 131, 136, 120, 124, 124, 125, 135, 122, 122, 118, 135, 121, 124, 132, 111, 116, 128, 125, 122, 119, 106, 138, 126, 124, 116, 116, 109, 115, 115, 128, 124, 115, 121, 123, 124, 116, 120, 112, 110, 116, 114, 119, 130, 131, 141, 149, 149, 140, 138, 122, 140, 147, 145, 147, 143, 141, 140, 125, 141, 126, 108, 116, 120, 125, 116, 116, 117, 112, 79, 67, 78, 81, 61, 58, 49, 58, 79, 88, 83, 83, 89, 85, 82, 76, 77, 72, 54, 49, 45, 48, 38, 39, 60, 79, 96, 100, 101, 101, 94, 95, 108, 100, 103, 103, 92, 102, 100, 108, 100, 99, 96, 93, 84, 97, 112, 96, 100, 99, 105, 105, 93, 101, 98, 106, 106, 99, 93, 101, 99, 99, 92, 99, 104, 108, 117, 122, 120, 124, 134, 124, 118, 127, 140, 132, 135, 128, 131, 120, 121, 126, 135, 140, 138, 139, 144, 142, 136, 127, 117, 111, 112, 117, 125, 121, 118, 114, 109, 128, 121, 121, 124, 110, 118, 119, 121, 121, 133, 128, 133, 134, 138, 141, 145, 144, 139, 149, 161, 141, 142, 151, 134, 144, 148, 152, 150, 157, 150, 154, 157, 161, 136, 146, 145, 153, 157, 159, 151, 160, 158, 129, 176, 158, 158, 163, 157, 126, 140, 151, 134, 132, 143, 133, 131, 132, 141, 133, 131, 123, 128, 131, 140, 140, 142, 137, 139, 134, 137, 141, 142, 139, 139, 125, 98, 165, 135, 135, 127, 135, 137, 129, 147, 133, 139, 135, 133, 138, 136, 135, 126, 132, 136, 138, 133, 118, 136, 114, 126, 119, 120, 120, 111, 104, 119, 117, 121, 125, 123, 127, 129, 126, 122, 121, 114, 112, 121, 124, 130, 123, 115, 121, 121, 124, 123, 114, 107, 119, 114, 121, 130, 128, 143, 155, 140, 147, 134, 136, 138, 142, 136, 139, 151, 144, 140, 130, 123, 129, 117, 118, 120, 127, 118, 111, 110, 101, 84, 75, 86, 85, 67, 56, 42, 43, 73, 77, 65, 75, 86, 91, 85, 72, 78, 77, 63, 44, 44, 49, 47, 40, 56, 80, 83, 91, 98, 96, 87, 95, 101, 106, 105, 106, 98, 93, 89, 113, 99, 99, 96, 92, 94, 94, 105, 93, 87, 95, 99, 90, 92, 94, 91, 93, 82, 100, 91, 92, 87, 102, 88, 100, 106, 106, 115, 117, 124, 145, 122, 109, 114, 130, 134, 134, 136, 129, 126, 118, 125, 127, 128, 134, 137, 133, 138, 140, 140, 131, 122, 113, 111, 108, 114, 120, 121, 120, 107, 126, 103, 110, 125, 108, 117, 112, 123, 124, 126, 125, 125, 132, 132, 133, 144, 147, 144, 138, 145, 135, 163, 140, 134, 144, 154, 146, 145, 153, 145, 157, 151, 152, 148, 146, 151, 153, 154, 157, 160, 154, 158, 156, 150, 168, 158, 163, 160, 120, 137, 142, 134, 141, 140, 138, 130, 124, 136, 128, 149, 133, 136, 125, 131, 139, 140, 135, 144, 136, 129, 145, 130, 140, 135, 139, 101, 136, 132, 131, 124, 126, 129, 144, 135, 139, 126, 137, 128, 131, 125, 122, 127, 123, 124, 129, 126, 123, 133, 124, 128, 122, 123, 118, 111, 120, 115, 128, 116, 120, 127, 128, 121, 117, 118, 123, 117, 117, 117, 126, 122, 121, 118, 125, 125, 122, 114, 109, 117, 112, 105, 138, 133, 133, 144, 161, 150, 154, 147, 144, 141, 146, 141, 118, 146, 144, 142, 133, 123, 121, 137, 116, 109, 116, 107, 110, 113, 104, 98, 96, 74, 74, 73, 67, 45, 44, 49, 60, 65, 65, 70, 73, 87, 87, 87, 79, 68, 55, 40, 45, 45, 42, 54, 59, 85, 98, 99, 102, 100, 97, 99, 107, 89, 123, 107, 95, 97, 99, 93, 94, 97, 88, 89, 93, 101, 85, 86, 91, 84, 101, 91, 89, 97, 93, 91, 90, 92, 78, 94, 93, 95, 100, 102, 110, 113, 115, 108, 131, 119, 114, 126, 122, 127, 142, 134, 128, 123, 126, 126, 127, 121, 119, 125, 127, 129, 133, 134, 138, 131, 126, 117, 122, 109, 118, 120, 117, 111, 110, 109, 108, 106, 107, 117, 104, 114, 123, 119, 131, 127, 134, 120, 137, 145, 131, 149, 138, 142, 130, 153, 129, 141, 151, 148, 149, 143, 145, 148, 153, 159, 156, 153, 151, 153, 153, 148, 152, 156, 153, 156, 154, 160, 169, 164, 158, 151, 129, 141, 126, 135, 134, 131, 134, 131, 132, 123, 119, 154, 156, 128, 144, 140, 136, 137, 119, 139, 133, 137, 147, 141, 141, 134, 136, 131, 138, 128, 131, 124, 129, 130, 137, 133, 138, 129, 135, 138, 126, 152, 119, 136, 145, 126, 126, 137, 124, 123, 115, 125, 131, 127, 119, 119, 125, 115, 120, 122, 116, 115, 105, 138, 121, 114, 111, 110, 117, 118, 123, 118, 126, 121, 116, 127, 135, 116, 115, 118, 112, 115, 129, 130, 130, 140, 147, 141, 166, 157, 145, 148, 144, 152, 145, 137, 138, 128, 132, 126, 123, 129, 120, 117, 120, 117, 107, 114, 96, 103, 98, 83, 65, 65, 58, 49, 45, 39, 53, 55, 49, 60, 76, 87, 90, 81, 80, 68, 52, 42, 58, 45, 46, 47, 55, 65, 88, 88, 100, 107, 89, 99, 112, 105, 108, 108, 101, 83, 88, 94, 85, 80, 82, 91, 94, 102, 95, 91, 95, 95, 92, 91, 89, 94, 91, 86, 96, 93, 94, 94, 84, 86, 89, 80, 106, 113, 102, 119, 119, 111, 151, 127, 127, 129, 128, 136, 121, 120, 124, 126, 133, 127, 126, 103, 126, 135, 120, 128, 136, 136, 121, 118, 127, 124, 116, 117, 116, 115, 118, 110, 118, 102, 111, 115, 109, 116, 123, 120, 125, 138, 132, 138, 135, 136, 137, 136, 141, 132, 147, 150, 139, 145, 149, 145, 142, 152, 148, 149, 151, 157, 150, 152, 155, 147, 158, 149, 149, 151, 130, 171, 148, 158, 157, 148, 156, 163, 137, 134, 131, 125, 126, 121, 124, 134, 123, 135, 116, 138, 135, 127, 150, 142, 135, 124, 143, 141, 131, 139, 141, 138, 139, 133, 133, 131, 135, 133, 121, 105, 130, 132, 136, 137, 133, 126, 127, 138, 128, 131, 126, 131, 138, 131, 131, 138, 135, 129, 130, 120, 122, 122, 121, 120, 120, 120, 120, 102, 110, 117, 108, 114, 117, 107, 117, 115, 137, 122, 124, 114, 125, 122, 122, 110, 129, 123, 127, 120, 120, 115, 123, 137, 140, 122, 139, 144, 155, 157, 156, 156, 152, 149, 146, 132, 146, 128, 127, 132, 122, 125, 118, 115, 120, 126, 114, 110, 111, 107, 97, 85, 65, 54, 48, 49, 46, 37, 34, 42, 53, 59, 64, 84, 89, 92, 88, 79, 55, 52, 58, 54, 51, 48, 47, 57, 75, 80, 91, 107, 95, 96, 106, 109, 105, 94, 91, 85, 86, 90, 78, 68, 83, 96, 93, 102, 95, 86, 98, 92, 93, 93, 86, 84, 86, 97, 93, 86, 101, 106, 90, 90, 93, 93, 112, 107, 98, 111, 100, 84, 140, 119, 128, 121, 132, 133, 124, 127, 124, 128, 126, 124, 123, 110, 127, 131, 117, 120, 127, 134, 110, 112, 136, 130, 120, 107, 112, 91, 105, 110, 110, 104, 102, 105, 123, 124, 125, 123, 127, 130, 134, 132, 141, 139, 133, 138, 139, 129, 148, 145, 143, 143, 146, 145, 144, 149, 147, 148, 145, 140, 146, 142, 158, 145, 146, 147, 145, 149, 140, 156, 154, 158, 143, 150, 152, 153, 128, 129, 134, 130, 122, 126, 120, 122, 138, 143, 137, 139, 135, 140, 139, 135, 137, 137, 136, 143, 136, 142, 137, 134, 139, 137, 134, 139, 133, 121, 124, 129, 122, 146, 129, 134, 112, 144, 147, 133, 131, 137, 137, 138, 135, 132, 133, 134, 130, 111, 145, 123, 121, 106, 116, 117, 119, 126, 120, 111, 115, 102, 112, 89, 118, 119, 117, 112, 130, 121, 128, 134, 125, 114, 119, 124, 128, 122, 117, 128, 123, 128, 123, 126, 141, 137, 121, 161, 158, 157, 161, 151, 146, 153, 141, 143, 137, 114, 121, 120, 129, 124, 112, 120, 120, 121, 120, 113, 112, 105, 95, 86, 67, 53, 54, 47, 44, 31, 19, 29, 43, 50, 56, 72, 83, 101, 86, 85, 70, 53, 50, 57, 47, 51, 53, 56, 60, 70, 83, 99, 89, 88, 99, 98, 105, 93, 83, 74, 94, 97, 88, 83, 97, 98, 97, 109, 101, 96, 88, 98, 93, 88, 89, 89, 94, 94, 93, 88, 97, 95, 91, 86, 100, 88, 119, 118, 115, 102, 101, 123, 127, 127, 121, 121, 134, 130, 118, 132, 121, 125, 122, 119, 131, 135, 120, 119, 126, 121, 120, 121, 115, 100, 109, 108, 100, 99, 111, 106, 106, 104, 107, 99, 103, 105, 124, 123, 136, 120, 132, 130, 128, 135, 132, 136, 135, 142, 139, 142, 141, 146, 148, 145, 141, 143, 147, 146, 149, 142, 146, 148, 144, 148, 146, 144, 142, 145, 145, 139, 144, 143, 149, 144, 148, 153, 149, 158, 131, 133, 129, 136, 128, 127, 135, 125, 135, 136, 142, 133, 142, 139, 141, 145, 139, 132, 140, 137, 137, 135, 141, 141, 134, 140, 141, 134, 136, 133, 124, 129, 135, 136, 137, 129, 124, 136, 132, 129, 136, 147, 126, 137, 135, 132, 126, 129, 132, 119, 134, 124, 124, 105, 114, 113, 113, 120, 117, 134, 121, 76, 108, 147, 141, 116, 120, 125, 125, 120, 129, 119, 112, 113, 119, 124, 117, 116, 119, 121, 118, 123, 127, 119, 130, 128, 139, 151, 165, 168, 161, 157, 161, 141, 138, 140, 134, 134, 127, 126, 127, 121, 116, 126, 119, 119, 118, 115, 110, 108, 103, 95, 70, 51, 50, 42, 29, 24, 19, 25, 32, 39, 50, 59, 70, 97, 94, 89, 68, 58, 59, 50, 32, 52, 66, 47, 53, 67, 83, 89, 85, 98, 99, 90, 95, 90, 93, 84, 91, 99, 93, 90, 101, 101, 94, 103, 109, 109, 85, 95, 84, 92, 90, 96, 91, 91, 92, 87, 95, 84, 96, 92, 100, 100, 114, 111, 107, 116, 124, 125, 125, 127, 131, 123, 123, 122, 125, 132, 119, 125, 122, 124, 136, 127, 123, 121, 123, 117, 127, 117, 121, 106, 107, 104, 102, 104, 107, 105, 110, 110, 108, 105, 110, 111, 125, 103, 133, 128, 127, 111, 122, 123, 127, 138, 137, 138, 140, 149, 139, 145, 145, 147, 144, 152, 149, 148, 147, 152, 131, 147, 148, 147, 146, 135, 122, 139, 126, 136, 160, 138, 138, 138, 140, 155, 145, 149, 138, 139, 129, 140, 134, 127, 138, 136, 138, 137, 138, 134, 141, 140, 136, 144, 141, 137, 136, 132, 124, 146, 142, 137, 137, 140, 143, 132, 135, 144, 132, 138, 136, 135, 145, 136, 129, 133, 125, 126, 131, 135, 127, 138, 129, 131, 122, 133, 128, 141, 121, 128, 125, 111, 120, 116, 120, 122, 116, 128, 122, 80, 99, 142, 137, 121, 123, 110, 132, 130, 118, 99, 106, 140, 136, 134, 117, 130, 122, 113, 113, 121, 109, 122, 132, 118, 149, 136, 153, 169, 157, 152, 170, 155, 139, 131, 134, 127, 121, 123, 122, 121, 123, 122, 118, 117, 126, 113, 117, 112, 116, 106, 82, 51, 41, 31, 20, 22, 16, 16, 25, 34, 43, 59, 70, 66, 104, 83, 83, 73, 53, 53, 41, 47, 53, 38, 51, 62, 74, 85, 77, 103, 85, 86, 89, 92, 92, 95, 92, 88, 95, 94, 94, 84, 92, 101, 87, 102, 92, 93, 81, 94, 87, 86, 81, 95, 83, 83, 86, 96, 88, 65, 97, 107, 111, 102, 116, 121, 133, 123, 125, 130, 126, 121, 120, 115, 115, 131, 128, 126, 125, 129, 124, 111, 108, 119, 99, 120, 122, 122, 127, 134, 119, 113, 95, 100, 115, 103, 109, 107, 111, 118, 114, 109, 123, 121, 121, 118, 118, 123, 134, 131, 140, 136, 136, 140, 133, 139, 141, 142, 149, 147, 152, 145, 146, 146, 129, 160, 146, 141, 148, 141, 138, 133, 107, 124, 116, 125, 159, 137, 133, 131, 152, 143, 147, 153, 139, 140, 133, 127, 135, 132, 131, 128, 157, 140, 134, 134, 136, 140, 144, 139, 132, 134, 138, 127, 134, 136, 134, 142, 140, 134, 137, 135, 133, 134, 137, 137, 134, 131, 130, 139, 140, 132, 138, 137, 127, 134, 127, 141, 135, 118, 136, 125, 137, 129, 101, 135, 118, 131, 120, 119, 121, 119, 119, 119, 122, 118, 107, 119, 113, 110, 120, 127, 125, 134, 104, 80, 112, 159, 182, 125, 107, 132, 120, 121, 109, 116, 101, 137, 141, 122, 146, 151, 154, 163, 167, 155, 156, 153, 140, 128, 118, 114, 111, 126, 128, 122, 119, 127, 132, 126, 124, 119, 118, 106, 105, 108, 81, 56, 37, 19, 13, 5, 11, 7, 2, 19, 38, 69, 74, 65, 88, 80, 80, 80, 63, 64, 50, 47, 49, 53, 49, 49, 56, 86, 88, 91, 77, 86, 88, 87, 92, 93, 87, 76, 94, 94, 93, 76, 102, 97, 99, 94, 97, 92, 86, 89, 92, 79, 92, 88, 83, 81, 87, 91, 80, 92, 109, 99, 99, 114, 127, 124, 122, 124, 117, 135, 123, 127, 127, 111, 122, 131, 130, 121, 104, 117, 126, 119, 115, 108, 85, 109, 128, 132, 136, 133, 115, 98, 115, 105, 109, 110, 111, 116, 106, 129, 137, 115, 124, 116, 121, 148, 118, 125, 131, 131, 139, 134, 126, 135, 146, 137, 133, 142, 141, 145, 143, 150, 141, 150, 143, 140, 137, 138, 139, 132, 132, 128, 120, 119, 119, 128, 149, 137, 141, 138, 144, 147, 148, 151, 124, 132, 133, 133, 129, 138, 134, 135, 149, 138, 137, 142, 134, 141, 138, 137, 132, 135, 138, 132, 131, 137, 129, 114, 139, 141, 139, 131, 139, 128, 139, 129, 121, 130, 135, 133, 131, 134, 127, 146, 139, 134, 128, 121, 146, 129, 131, 138, 134, 116, 130, 119, 125, 125, 133, 117, 110, 118, 110, 122, 122, 133, 123, 127, 121, 112, 113, 121, 126, 128, 78, 74, 117, 157, 178, 129, 119, 124, 121, 123, 101, 119, 118, 121, 116, 121, 143, 150, 155, 175, 170, 164, 158, 143, 145, 134, 118, 100, 110, 121, 127, 128, 116, 126, 139, 130, 126, 127, 110, 108, 99, 100, 77, 53, 33, 23, 17, 9, 6, 9, 6, 11, 3, 45, 71, 72, 76, 85, 75, 71, 70, 58, 41, 52, 50, 44, 44, 50, 58, 80, 98, 80, 67, 83, 93, 97, 95, 99, 90, 87, 96, 99, 86, 92, 94, 97, 88, 95, 97, 89, 83, 81, 94, 97, 92, 84, 103, 99, 88, 91, 87, 91, 95, 98, 81, 106, 130, 128, 119, 120, 98, 138, 129, 125, 130, 119, 121, 115, 129, 117, 107, 115, 127, 124, 127, 113, 90, 105, 119, 137, 137, 119, 109, 92, 113, 108, 105, 112, 112, 121, 89, 128, 167, 119, 122, 119, 116, 118, 123, 127, 132, 133, 130, 131, 153, 137, 147, 144, 133, 140, 135, 139, 142, 144, 145, 148, 143, 137, 143, 143, 141, 136, 134, 135, 126, 104, 125, 162, 143, 127, 124, 130, 151, 148, 154, 146, 131, 134, 137, 136, 138, 137, 137, 139, 135, 136, 138, 141, 141, 135, 147, 143, 142, 141, 135, 127, 143, 135, 137, 127, 134, 137, 139, 133, 139, 134, 135, 135, 133, 135, 108, 159, 129, 132, 131, 132, 130, 133, 143, 126, 134, 126, 132, 135, 137, 141, 123, 127, 126, 120, 126, 126, 112, 118, 108, 116, 116, 132, 125, 124, 123, 113, 124, 120, 123, 128, 94, 77, 122, 139, 153, 118, 118, 122, 121, 120, 116, 110, 122, 124, 123, 125, 146, 156, 157, 169, 175, 171, 165, 148, 136, 128, 115, 95, 90, 112, 131, 133, 121, 122, 138, 128, 131, 133, 120, 108, 97, 79, 70, 56, 30, 19, 13, 4, 0, 4, 10, 7, 14, 34, 58, 66, 70, 75, 68, 59, 63, 59, 47, 48, 46, 50, 48, 48, 56, 78, 82, 74, 67, 75, 92, 92, 100, 100, 99, 96, 104, 100, 93, 97, 97, 93, 83, 87, 92, 96, 88, 88, 96, 96, 80, 73, 113, 113, 86, 99, 92, 81, 94, 96, 91, 115, 111, 117, 122, 120, 122, 128, 130, 110, 120, 113, 115, 113, 109, 110, 106, 98, 102, 114, 129, 119, 97, 112, 128, 135, 118, 110, 108, 103, 116, 122, 117, 109, 119, 119, 88, 113, 139, 113, 120, 121, 118, 116, 120, 131, 130, 128, 140, 132, 137, 132, 132, 137, 155, 142, 142, 147, 144, 138, 140, 143, 136, 142, 147, 139, 139, 139, 137, 141, 136, 143, 130, 137, 138, 134, 132, 144, 148, 147, 151, 157, 136, 132, 140, 138, 135, 141, 137, 135, 136, 131, 137, 137, 143, 140, 140, 142, 138, 134, 135, 136, 130, 137, 141, 134, 136, 137, 134, 137, 139, 133, 137, 136, 133, 135, 122, 138, 131, 130, 135, 134, 128, 134, 128, 137, 119, 118, 129, 135, 132, 135, 126, 126, 134, 114, 124, 115, 118, 117, 110, 121, 116, 107, 112, 124, 123, 121, 116, 132, 128, 128, 115, 98, 109, 134, 125, 110, 115, 124, 124, 118, 116, 124, 113, 118, 134, 114, 137, 154, 151, 170, 179, 176, 163, 160, 134, 121, 98, 97, 80, 97, 126, 119, 106, 129, 138, 135, 139, 135, 129, 108, 101, 81, 57, 39, 26, 14, 4, 0, 0, 3, 13, 7, 8, 25, 44, 54, 66, 60, 60, 64, 54, 43, 42, 44, 36, 37, 49, 55, 58, 69, 78, 77, 75, 80, 86, 94, 95, 101, 104, 96, 98, 103, 93, 100, 104, 95, 87, 89, 88, 83, 101, 99, 101, 101, 78, 74, 107, 114, 97, 90, 83, 83, 93, 104, 98, 112, 121, 116, 114, 128, 120, 119, 108, 113, 112, 104, 105, 110, 109, 104, 86, 84, 106, 119, 131, 115, 113, 107, 122, 124, 112, 109, 112, 108, 110, 124, 116, 110, 122, 117, 117, 114, 119, 115, 123, 126, 120, 116, 128, 130, 129, 125, 137, 130, 131, 135, 132, 137, 148, 140, 142, 139, 138, 138, 148, 117, 169, 136, 140, 137, 139, 139, 138, 136, 143, 139, 140, 142, 143, 147, 149, 151, 154, 158, 152, 147, 135, 134, 135, 136, 129, 139, 132, 140, 128, 131, 139, 140, 139, 140, 142, 145, 138, 130, 128, 137, 137, 136, 121, 138, 134, 131, 135, 130, 137, 139, 138, 131, 132, 139, 141, 127, 137, 137, 133, 130, 137, 137, 130, 133, 121, 128, 127, 127, 133, 127, 132, 136, 131, 125, 119, 123, 120, 123, 116, 116, 113, 110, 115, 108, 121, 122, 115, 128, 125, 123, 117, 122, 118, 124, 116, 123, 120, 125, 126, 121, 113, 127, 122, 104, 125, 136, 132, 140, 161, 170, 179, 172, 161, 155, 134, 120, 113, 117, 91, 97, 115, 115, 119, 116, 139, 160, 152, 146, 135, 124, 117, 89, 64, 45, 19, 18, 6, 0, 0, 0, 3, 15, 14, 25, 37, 48, 50, 50, 48, 50, 50, 48, 44, 37, 32, 38, 32, 40, 54, 64, 73, 70, 76, 87, 87, 99, 102, 99, 107, 100, 103, 99, 95, 95, 95, 98, 91, 98, 92, 95, 95, 98, 98, 101, 90, 96, 101, 101, 102, 98, 97, 97, 100, 87, 91, 117, 148, 145, 117, 119, 121, 120, 115, 119, 120, 107, 89, 108, 116, 98, 77, 81, 91, 109, 119, 118, 124, 98, 121, 121, 115, 114, 117, 118, 117, 118, 111, 110, 122, 121, 120, 108, 122, 122, 112, 125, 123, 117, 110, 121, 126, 115, 144, 128, 133, 138, 128, 135, 133, 128, 136, 126, 140, 144, 144, 126, 147, 137, 134, 140, 129, 138, 132, 133, 142, 148, 140, 145, 144, 149, 159, 155, 153, 157, 152, 161, 132, 149, 139, 134, 136, 136, 125, 148, 137, 137, 137, 137, 135, 139, 137, 126, 139, 131, 118, 125, 142, 131, 76, 138, 170, 120, 132, 142, 133, 138, 133, 131, 124, 129, 136, 127, 135, 126, 116, 134, 131, 134, 128, 126, 132, 130, 125, 130, 128, 137, 132, 128, 126, 122, 132, 117, 118, 116, 120, 110, 137, 117, 127, 125, 118, 118, 121, 128, 116, 121, 126, 124, 122, 118, 121, 114, 126, 123, 103, 133, 100, 128, 116, 108, 116, 117, 119, 140, 150, 167, 169, 172, 170, 156, 135, 122, 112, 118, 109, 105, 106, 103, 111, 101, 147, 164, 165, 148, 142, 137, 116, 102, 63, 48, 26, 11, 1, 0, 0, 0, 0, 16, 11, 17, 33, 38, 43, 43, 36, 34, 35, 41, 36, 38, 29, 26, 26, 33, 48, 52, 65, 72, 74, 78, 85, 100, 88, 111, 108, 102, 99, 107, 102, 96, 90, 100, 90, 88, 86, 99, 94, 97, 100, 95, 85, 101, 98, 96, 101, 103, 105, 104, 93, 80, 80, 114, 146, 153, 125, 111, 115, 117, 109, 111, 117, 109, 99, 107, 102, 85, 64, 96, 83, 98, 101, 111, 134, 118, 112, 124, 118, 116, 116, 128, 115, 116, 125, 110, 127, 116, 122, 112, 128, 124, 115, 114, 121, 126, 122, 118, 117, 108, 136, 125, 128, 129, 133, 134, 137, 129, 131, 140, 141, 150, 142, 138, 127, 148, 143, 139, 136, 144, 131, 132, 129, 140, 140, 138, 152, 150, 150, 151, 160, 150, 154, 157, 123, 139, 131, 138, 139, 134, 135, 123, 149, 141, 139, 133, 120, 126, 126, 129, 135, 138, 126, 122, 130, 136, 108, 114, 132, 123, 137, 137, 130, 129, 131, 126, 139, 131, 135, 123, 123, 128, 110, 130, 126, 136, 125, 131, 128, 123, 128, 118, 130, 117, 127, 119, 125, 119, 118, 123, 113, 122, 124, 112, 122, 123, 114, 120, 125, 109, 126, 135, 123, 128, 124, 127, 127, 119, 126, 123, 118, 130, 116, 108, 115, 117, 105, 117, 142, 119, 118, 140, 139, 161, 164, 161, 173, 152, 132, 120, 101, 118, 109, 100, 105, 110, 91, 80, 127, 156, 167, 163, 154, 137, 123, 95, 67, 50, 29, 5, 1, 6, 0, 1, 0, 10, 5, 11, 20, 32, 58, 54, 39, 30, 33, 32, 28, 30, 20, 18, 23, 29, 38, 44, 56, 65, 71, 75, 81, 92, 95, 104, 105, 106, 96, 97, 102, 97, 92, 97, 98, 102, 90, 85, 83, 101, 90, 96, 110, 106, 99, 104, 105, 108, 106, 103, 112, 78, 82, 113, 134, 143, 108, 113, 110, 118, 108, 110, 110, 111, 105, 108, 80, 73, 77, 110, 108, 108, 98, 106, 130, 112, 113, 118, 120, 117, 118, 117, 120, 116, 124, 100, 121, 97, 124, 111, 121, 116, 112, 109, 101, 126, 124, 115, 109, 122, 130, 126, 124, 132, 127, 133, 137, 139, 143, 140, 143, 136, 144, 135, 137, 138, 141, 131, 127, 132, 137, 128, 132, 141, 140, 140, 150, 155, 157, 154, 158, 154, 157, 161, 146, 137, 127, 140, 140, 138, 135, 133, 139, 136, 137, 122, 115, 126, 125, 127, 124, 130, 125, 133, 125, 125, 134, 124, 139, 131, 132, 135, 142, 116, 130, 135, 130, 126, 127, 125, 125, 125, 126, 126, 126, 121, 117, 126, 107, 102, 153, 131, 115, 127, 126, 119, 120, 113, 120, 117, 120, 107, 119, 121, 125, 123, 115, 124, 116, 127, 113, 126, 120, 129, 118, 122, 116, 127, 125, 119, 121, 125, 124, 119, 125, 118, 110, 112, 129, 121, 122, 139, 144, 154, 165, 171, 165, 145, 138, 126, 111, 114, 99, 83, 92, 109, 107, 79, 112, 160, 167, 162, 172, 145, 139, 108, 84, 58, 18, 11, 0, 0, 0, 0, 0, 4, 7, 4, 7, 26, 74, 77, 30, 20, 29, 32, 26, 20, 20, 15, 18, 27, 39, 36, 46, 56, 66, 84, 83, 94, 99, 97, 104, 96, 97, 100, 104, 99, 95, 91, 99, 105, 98, 92, 88, 93, 91, 101, 111, 106, 108, 99, 109, 95, 84, 101, 109, 101, 80, 106, 119, 116, 106, 118, 126, 117, 116, 114, 110, 111, 93, 99, 80, 69, 85, 104, 117, 105, 104, 108, 120, 113, 108, 114, 117, 124, 118, 114, 118, 114, 119, 108, 114, 107, 117, 116, 109, 109, 106, 144, 114, 130, 124, 110, 122, 115, 125, 123, 113, 143, 137, 133, 129, 137, 138, 135, 134, 129, 144, 135, 136, 124, 131, 136, 125, 131, 137, 129, 128, 141, 140, 150, 145, 145, 152, 160, 157, 144, 149, 176, 135, 140, 137, 137, 140, 135, 135, 130, 131, 129, 135, 126, 127, 128, 131, 133, 125, 131, 132, 125, 130, 139, 134, 138, 138, 128, 137, 139, 128, 134, 134, 127, 126, 126, 132, 120, 107, 103, 125, 123, 122, 118, 125, 123, 100, 89, 140, 154, 117, 124, 116, 114, 121, 117, 112, 115, 120, 127, 108, 112, 119, 125, 113, 124, 116, 117, 122, 125, 126, 125, 123, 123, 105, 123, 120, 123, 122, 124, 127, 125, 121, 124, 108, 110, 115, 117, 112, 132, 144, 150, 160, 170, 179, 149, 133, 125, 110, 104, 78, 55, 76, 115, 158, 139, 132, 163, 168, 173, 162, 164, 161, 107, 88, 63, 21, 11, 0, 0, 0, 0, 0, 0, 5, 0, 1, 14, 83, 91, 27, 13, 31, 50, 36, 18, 17, 19, 16, 18, 17, 26, 34, 42, 55, 69, 72, 89, 98, 97, 96, 94, 97, 98, 102, 99, 106, 98, 102, 103, 94, 97, 97, 93, 102, 101, 106, 101, 109, 119, 107, 101, 106, 115, 115, 106, 101, 107, 111, 112, 106, 116, 125, 117, 112, 103, 112, 115, 104, 100, 82, 66, 91, 100, 103, 86, 93, 123, 117, 122, 112, 117, 114, 125, 123, 117, 109, 116, 104, 107, 115, 110, 117, 109, 109, 116, 90, 116, 110, 154, 127, 113, 108, 124, 122, 116, 104, 147, 148, 116, 125, 135, 136, 132, 122, 135, 136, 137, 128, 125, 133, 133, 135, 127, 133, 137, 136, 149, 152, 153, 154, 146, 166, 160, 155, 140, 152, 172, 145, 145, 130, 138, 137, 140, 127, 129, 125, 128, 143, 129, 127, 128, 128, 129, 132, 134, 131, 134, 120, 127, 149, 137, 131, 135, 133, 136, 127, 129, 126, 142, 123, 129, 130, 119, 98, 116, 125, 127, 128, 115, 117, 119, 112, 96, 121, 123, 116, 127, 111, 113, 115, 113, 96, 104, 109, 143, 109, 116, 124, 119, 125, 126, 124, 120, 125, 121, 124, 117, 120, 121, 127, 119, 117, 116, 119, 123, 118, 106, 103, 124, 140, 125, 109, 121, 105, 122, 134, 135, 152, 168, 184, 157, 128, 126, 121, 100, 52, 33, 63, 104, 172, 179, 129, 143, 161, 171, 165, 164, 158, 120, 84, 53, 31, 12, 1, 0, 6, 14, 0, 4, 4, 0, 0, 17, 71, 68, 12, 3, 17, 65, 55, 22, 13, 14, 6, 12, 7, 11, 16, 26, 54, 53, 74, 87, 88, 96, 96, 99, 94, 99, 98, 104, 99, 102, 96, 102, 99, 99, 98, 95, 96, 104, 103, 103, 107, 111, 92, 99, 106, 114, 110, 104, 106, 111, 117, 117, 117, 116, 126, 119, 103, 105, 105, 119, 109, 98, 86, 79, 97, 91, 94, 81, 99, 127, 122, 120, 114, 110, 114, 120, 118, 123, 117, 108, 109, 117, 109, 109, 125, 109, 103, 115, 110, 116, 113, 124, 122, 124, 99, 106, 108, 122, 97, 135, 127, 126, 130, 126, 135, 132, 127, 131, 128, 127, 125, 123, 116, 127, 132, 133, 146, 147, 146, 151, 156, 161, 155, 154, 157, 156, 158, 152, 156, 157, 136, 138, 134, 136, 132, 134, 128, 129, 132, 126, 128, 135, 137, 136, 107, 127, 134, 124, 129, 131, 126, 121, 133, 128, 128, 136, 126, 127, 138, 131, 113, 128, 115, 122, 120, 118, 111, 122, 124, 117, 120, 118, 113, 112, 118, 115, 107, 111, 115, 118, 116, 113, 84, 91, 88, 94, 83, 117, 114, 126, 124, 122, 128, 125, 123, 128, 120, 118, 116, 125, 113, 117, 124, 116, 131, 131, 110, 119, 132, 85, 88, 119, 167, 156, 110, 110, 107, 106, 134, 131, 143, 175, 178, 174, 139, 119, 114, 92, 49, 32, 45, 88, 157, 173, 127, 142, 160, 176, 176, 171, 165, 130, 88, 48, 32, 7, 10, 3, 9, 27, 11, 6, 16, 4, 0, 14, 39, 34, 10, 0, 7, 56, 49, 14, 16, 7, 3, 11, 2, 3, 16, 29, 54, 54, 75, 90, 88, 94, 95, 96, 99, 98, 99, 103, 99, 104, 97, 103, 106, 108, 102, 103, 105, 105, 102, 107, 110, 103, 95, 99, 108, 110, 109, 110, 106, 113, 112, 124, 120, 115, 118, 105, 109, 108, 110, 125, 114, 96, 97, 86, 90, 97, 95, 105, 107, 121, 121, 124, 118, 109, 121, 117, 117, 118, 115, 107, 98, 111, 115, 107, 119, 108, 108, 108, 111, 112, 128, 110, 115, 117, 113, 113, 97, 123, 119, 125, 123, 119, 127, 136, 131, 133, 137, 134, 136, 120, 114, 130, 134, 139, 143, 148, 142, 153, 148, 149, 152, 155, 150, 150, 155, 155, 160, 155, 147, 157, 138, 136, 138, 137, 133, 129, 131, 123, 137, 135, 139, 138, 137, 131, 136, 129, 126, 127, 135, 126, 128, 123, 130, 124, 133, 122, 132, 114, 142, 121, 124, 121, 112, 109, 106, 113, 106, 109, 112, 119, 109, 107, 115, 106, 112, 114, 115, 90, 106, 102, 80, 84, 119, 70, 70, 100, 93, 103, 107, 116, 116, 122, 122, 122, 125, 123, 126, 125, 119, 129, 107, 121, 118, 105, 128, 119, 111, 121, 114, 83, 77, 117, 153, 162, 112, 117, 110, 101, 127, 136, 135, 164, 171, 163, 141, 117, 113, 93, 57, 31, 47, 83, 123, 126, 100, 128, 161, 168, 170, 176, 163, 119, 87, 77, 33, 10, 5, 15, 4, 18, 34, 13, 14, 14, 15, 29, 37, 19, 6, 0, 9, 30, 35, 24, 10, 2, 11, 32, 11, 9, 14, 31, 51, 63, 77, 78, 86, 107, 91, 90, 94, 102, 104, 106, 99, 101, 102, 101, 100, 100, 110, 105, 104, 99, 98, 107, 109, 102, 93, 99, 108, 110, 107, 107, 111, 111, 104, 118, 124, 115, 126, 111, 107, 111, 119, 117, 122, 85, 120, 98, 103, 106, 94, 108, 117, 116, 121, 117, 116, 113, 122, 119, 112, 123, 120, 103, 119, 111, 112, 110, 111, 101, 108, 117, 121, 114, 127, 107, 126, 104, 106, 94, 99, 107, 125, 119, 127, 130, 130, 132, 129, 136, 130, 131, 126, 116, 125, 140, 137, 148, 146, 149, 147, 150, 150, 149, 155, 161, 150, 159, 152, 146, 156, 150, 159, 159, 138, 135, 138, 132, 132, 134, 137, 125, 130, 133, 138, 127, 134, 131, 135, 135, 131, 126, 118, 130, 124, 120, 124, 128, 121, 128, 129, 125, 128, 117, 133, 108, 94, 98, 101, 108, 88, 111, 122, 97, 113, 98, 100, 106, 85, 108, 108, 100, 113, 104, 68, 71, 98, 91, 88, 68, 87, 116, 104, 118, 125, 116, 119, 116, 126, 122, 118, 110, 123, 131, 108, 111, 111, 117, 128, 101, 116, 141, 126, 88, 85, 114, 144, 140, 99, 113, 113, 106, 113, 140, 131, 138, 167, 157, 138, 108, 97, 93, 94, 74, 54, 73, 96, 81, 91, 134, 158, 169, 165, 161, 158, 117, 94, 74, 40, 12, 11, 30, 20, 21, 22, 19, 18, 15, 22, 41, 31, 18, 13, 12, 10, 13, 30, 33, 6, 1, 15, 39, 17, 2, 9, 23, 30, 54, 67, 62, 80, 119, 98, 104, 95, 94, 105, 98, 103, 99, 99, 98, 96, 101, 109, 98, 102, 103, 105, 106, 107, 104, 103, 94, 92, 134, 154, 121, 111, 112, 102, 116, 121, 127, 127, 111, 112, 116, 113, 120, 115, 92, 90, 78, 92, 101, 105, 116, 114, 106, 118, 113, 115, 120, 123, 109, 108, 120, 119, 124, 117, 115, 114, 108, 98, 124, 109, 112, 117, 109, 116, 105, 118, 117, 105, 101, 102, 130, 122, 124, 117, 127, 134, 135, 132, 133, 127, 133, 139, 136, 141, 138, 146, 149, 149, 149, 144, 149, 154, 149, 148, 160, 149, 153, 140, 149, 163, 155, 156, 160, 129, 138, 135, 120, 144, 137, 124, 128, 137, 119, 125, 138, 135, 135, 138, 130, 131, 126, 115, 123, 134, 117, 126, 129, 125, 120, 124, 127, 122, 106, 121, 98, 73, 95, 107, 106, 91, 103, 111, 98, 115, 94, 100, 99, 92, 107, 110, 106, 112, 101, 79, 81, 116, 102, 84, 99, 101, 109, 121, 104, 113, 115, 102, 141, 119, 119, 117, 117, 118, 118, 111, 117, 118, 119, 124, 104, 114, 128, 124, 119, 102, 101, 118, 103, 106, 112, 111, 109, 111, 127, 129, 128, 147, 141, 122, 119, 93, 79, 115, 124, 95, 71, 90, 102, 86, 126, 160, 173, 168, 164, 144, 124, 103, 68, 46, 22, 21, 43, 21, 28, 19, 20, 16, 29, 18, 16, 16, 12, 19, 19, 10, 26, 36, 50, 26, 22, 25, 23, 11, 0, 2, 9, 29, 42, 67, 74, 79, 101, 98, 97, 102, 102, 102, 101, 95, 87, 103, 107, 101, 98, 112, 95, 94, 112, 105, 108, 112, 105, 95, 77, 81, 134, 170, 144, 107, 117, 117, 116, 118, 120, 123, 101, 93, 99, 117, 123, 117, 106, 86, 85, 91, 88, 102, 120, 117, 109, 111, 112, 108, 121, 111, 105, 112, 105, 115, 123, 110, 122, 120, 106, 110, 122, 111, 114, 115, 118, 114, 116, 114, 108, 124, 110, 123, 123, 129, 126, 127, 135, 133, 134, 141, 146, 128, 138, 129, 136, 148, 137, 145, 148, 152, 145, 148, 145, 151, 156, 150, 151, 153, 155, 157, 155, 146, 154, 150, 164, 129, 133, 135, 128, 138, 127, 132, 129, 132, 131, 138, 130, 131, 133, 127, 126, 131, 128, 125, 127, 132, 120, 123, 125, 110, 117, 124, 115, 115, 102, 112, 105, 99, 101, 105, 111, 100, 114, 107, 107, 104, 103, 92, 110, 98, 102, 102, 109, 106, 109, 82, 83, 133, 113, 85, 112, 99, 112, 110, 115, 115, 117, 116, 118, 105, 127, 118, 117, 118, 126, 116, 116, 118, 120, 126, 114, 116, 120, 106, 127, 107, 115, 109, 109, 97, 115, 110, 106, 103, 125, 135, 129, 141, 135, 127, 115, 90, 65, 98, 109, 96, 67, 79, 136, 152, 134, 151, 169, 162, 164, 143, 117, 99, 75, 61, 41, 39, 37, 33, 30, 34, 39, 35, 47, 30, 25, 18, 10, 22, 17, 14, 13, 27, 42, 50, 58, 30, 1, 11, 1, 0, 3, 11, 28, 59, 79, 91, 94, 97, 83, 108, 110, 104, 109, 98, 88, 99, 104, 105, 107, 102, 103, 98, 102, 108, 100, 113, 110, 104, 83, 82, 115, 152, 122, 114, 116, 116, 116, 126, 123, 122, 106, 98, 99, 111, 138, 108, 99, 93, 92, 88, 93, 117, 117, 112, 116, 117, 113, 116, 121, 107, 116, 119, 111, 114, 121, 99, 126, 120, 113, 113, 118, 121, 114, 114, 118, 118, 121, 125, 120, 119, 118, 127, 131, 119, 127, 135, 133, 137, 136, 137, 139, 146, 137, 139, 141, 147, 143, 144, 147, 149, 151, 144, 139, 151, 155, 142, 159, 146, 150, 152, 152, 153, 160, 150, 157, 140, 137, 137, 140, 129, 126, 136, 137, 136, 132, 139, 126, 137, 119, 122, 123, 127, 129, 133, 133, 132, 138, 130, 129, 118, 126, 118, 113, 111, 108, 109, 103, 95, 109, 109, 116, 111, 125, 104, 94, 108, 99, 105, 102, 105, 108, 105, 96, 101, 81, 65, 92, 155, 139, 106, 111, 91, 131, 135, 107, 112, 114, 114, 114, 113, 119, 115, 116, 116, 118, 120, 115, 114, 118, 112, 121, 120, 116, 106, 111, 99, 113, 100, 112, 104, 103, 99, 108, 106, 120, 127, 109, 116, 137, 148, 142, 108, 85, 62, 84, 101, 84, 75, 144, 181, 159, 152, 169, 161, 155, 139, 128, 122, 87, 70, 62, 57, 50, 44, 34, 48, 66, 61, 47, 37, 27, 26, 11, 7, 1, 5, 10, 28, 42, 67, 61, 25, 5, 3, 0, 0, 0, 1, 13, 44, 76, 69, 89, 97, 83, 91, 91, 138, 153, 110, 89, 95, 100, 106, 114, 112, 107, 104, 102, 108, 109, 116, 117, 117, 101, 86, 104, 125, 105, 99, 117, 113, 118, 127, 112, 117, 108, 102, 88, 90, 126, 98, 96, 97, 98, 111, 105, 108, 116, 119, 119, 112, 114, 123, 117, 111, 114, 120, 118, 119, 118, 110, 114, 122, 114, 114, 125, 124, 114, 116, 119, 111, 117, 119, 126, 128, 121, 128, 124, 128, 128, 134, 123, 147, 144, 143, 147, 141, 150, 148, 144, 144, 136, 146, 145, 146, 145, 153, 148, 148, 153, 161, 159, 151, 154, 151, 157, 154, 153, 157, 164, 130, 132, 142, 132, 134, 132, 131, 135, 140, 124, 133, 128, 135, 117, 119, 118, 133, 132, 131, 133, 131, 130, 130, 127, 120, 122, 121, 118, 118, 121, 117, 114, 106, 113, 116, 108, 104, 95, 103, 85, 116, 95, 113, 103, 102, 103, 103, 101, 103, 104, 63, 104, 155, 133, 112, 115, 77, 125, 160, 117, 111, 118, 112, 119, 122, 117, 115, 112, 116, 125, 112, 112, 103, 117, 111, 115, 113, 116, 106, 111, 94, 118, 111, 109, 112, 98, 101, 90, 98, 115, 108, 75, 92, 126, 163, 164, 136, 98, 51, 61, 95, 105, 74, 150, 181, 163, 141, 155, 168, 164, 140, 121, 118, 93, 79, 67, 64, 59, 41, 41, 50, 66, 69, 58, 37, 32, 33, 7, 0, 13, 20, 14, 29, 50, 68, 45, 4, 3, 0, 0, 0, 16, 17, 14, 29, 68, 77, 88, 89, 88, 66, 66, 120, 167, 148, 96, 95, 95, 101, 99, 90, 103, 101, 104, 107, 114, 116, 110, 113, 124, 108, 108, 117, 106, 110, 112, 124, 119, 119, 124, 113, 99, 103, 104, 108, 110, 106, 101, 102, 105, 118, 110, 110, 121, 126, 120, 120, 120, 115, 116, 115, 114, 121, 115, 112, 118, 116, 110, 113, 110, 110, 119, 126, 110, 117, 122, 113, 112, 118, 113, 127, 124, 132, 122, 140, 126, 136, 134, 147, 133, 143, 145, 143, 147, 152, 151, 143, 147, 150, 143, 147, 149, 151, 149, 153, 154, 151, 156, 160, 152, 155, 155, 151, 155, 159, 152, 136, 139, 137, 135, 128, 133, 128, 131, 135, 133, 135, 135, 135, 131, 132, 130, 133, 131, 129, 122, 128, 134, 126, 125, 123, 127, 113, 120, 122, 120, 125, 116, 119, 105, 102, 118, 117, 109, 108, 110, 106, 104, 111, 98, 110, 99, 65, 88, 110, 137, 92, 83, 135, 95, 112, 108, 92, 116, 131, 107, 113, 105, 108, 108, 112, 111, 111, 107, 109, 116, 109, 114, 97, 109, 108, 114, 102, 119, 111, 110, 103, 114, 112, 106, 111, 104, 99, 70, 77, 96, 102, 68, 67, 111, 160, 161, 124, 98, 73, 62, 99, 93, 73, 109, 178, 154, 116, 131, 181, 180, 154, 121, 103, 93, 77, 66, 85, 68, 45, 42, 58, 72, 77, 60, 38, 26, 38, 14, 0, 15, 44, 15, 29, 50, 61, 52, 23, 6, 0, 0, 0, 21, 32, 13, 18, 51, 77, 88, 94, 98, 59, 49, 99, 142, 129, 99, 103, 91, 95, 104, 99, 105, 109, 100, 116, 103, 107, 111, 124, 121, 101, 105, 111, 111, 102, 100, 117, 112, 115, 115, 114, 112, 99, 104, 108, 81, 132, 99, 99, 112, 114, 122, 102, 119, 119, 117, 113, 112, 115, 116, 117, 116, 117, 117, 109, 116, 116, 115, 112, 114, 110, 117, 118, 118, 123, 115, 114, 115, 122, 129, 124, 129, 135, 126, 128, 136, 140, 136, 131, 154, 138, 149, 141, 150, 149, 152, 141, 149, 148, 144, 152, 153, 141, 161, 163, 151, 155, 155, 151, 157, 153, 155, 157, 142, 160, 146, 134, 136, 128, 138, 132, 133, 127, 133, 128, 134, 131, 128, 128, 131, 127, 132, 137, 126, 131, 124, 124, 129, 133, 129, 130, 130, 129, 119, 137, 125, 121, 120, 122, 111, 109, 110, 114, 104, 117, 114, 101, 106, 109, 116, 95, 88, 70, 79, 109, 104, 123, 111, 109, 105, 114, 117, 127, 97, 114, 114, 98, 114, 107, 110, 108, 114, 97, 118, 110, 109, 108, 103, 108, 107, 111, 111, 105, 109, 115, 112, 111, 107, 111, 101, 112, 112, 112, 97, 101, 97, 85, 83, 68, 81, 125, 132, 116, 94, 100, 95, 100, 96, 81, 89, 152, 137, 97, 96, 185, 188, 152, 123, 114, 83, 80, 72, 76, 76, 65, 56, 64, 75, 69, 55, 44, 48, 33, 7, 0, 20, 24, 6, 34, 42, 26, 51, 34, 23, 3, 0, 0, 19, 12, 1, 18, 31, 70, 92, 93, 109, 74, 53, 85, 119, 91, 91, 105, 105, 104, 106, 106, 103, 106, 109, 111, 111, 108, 104, 125, 115, 100, 106, 103, 111, 109, 94, 103, 111, 121, 109, 92, 135, 103, 109, 106, 97, 107, 93, 106, 115, 124, 121, 112, 102, 117, 117, 107, 116, 124, 102, 120, 118, 110, 118, 109, 111, 105, 135, 119, 110, 116, 119, 119, 119, 110, 117, 121, 117, 109, 119, 116, 127, 130, 134, 141, 136, 134, 140, 127, 145, 141, 147, 143, 145, 152, 149, 144, 146, 144, 140, 148, 151, 144, 153, 157, 152, 159, 157, 148, 153, 155, 154, 158, 158, 160, 155, 107, 153, 144, 131, 135, 138, 127, 119, 130, 132, 139, 128, 134, 133, 136, 128, 133, 119, 134, 129, 121, 133, 138, 134, 127, 107, 130, 132, 129, 125, 117, 127, 114, 119, 118, 114, 105, 117, 108, 109, 97, 105, 96, 100, 90, 85, 67, 85, 98, 77, 124, 94, 112, 104, 99, 122, 132, 107, 102, 80, 96, 108, 106, 104, 117, 111, 109, 103, 105, 95, 102, 109, 107, 111, 98, 106, 104, 101, 104, 103, 101, 118, 109, 112, 104, 123, 112, 102, 105, 108, 98, 105, 93, 90, 99, 97, 86, 106, 107, 88, 104, 115, 92, 122, 145, 136, 105, 94, 158, 168, 141, 124, 116, 83, 80, 85, 84, 76, 78, 70, 67, 73, 75, 68, 45, 45, 33, 18, 14, 42, 28, 13, 21, 34, 33, 31, 32, 9, 0, 0, 3, 4, 1, 3, 21, 30, 50, 92, 93, 96, 94, 86, 84, 108, 89, 101, 107, 99, 106, 107, 115, 115, 111, 108, 108, 104, 112, 113, 120, 112, 112, 106, 102, 112, 104, 113, 101, 121, 105, 95, 109, 126, 121, 114, 102, 105, 97, 103, 107, 119, 117, 126, 117, 103, 124, 117, 114, 110, 115, 119, 116, 110, 117, 120, 114, 117, 110, 117, 108, 115, 113, 108, 118, 115, 112, 121, 119, 124, 116, 124, 133, 126, 124, 134, 132, 140, 141, 135, 148, 139, 134, 144, 156, 149, 142, 152, 145, 150, 133, 141, 149, 149, 148, 156, 151, 159, 150, 153, 145, 161, 153, 152, 146, 151, 152, 147, 111, 127, 151, 129, 128, 131, 129, 118, 129, 128, 135, 116, 156, 123, 127, 143, 131, 124, 130, 140, 128, 133, 126, 132, 132, 100, 145, 125, 111, 119, 125, 123, 117, 118, 114, 107, 110, 99, 111, 99, 106, 100, 105, 101, 92, 87, 75, 77, 87, 108, 113, 109, 109, 114, 94, 115, 106, 102, 108, 82, 79, 89, 109, 101, 114, 107, 108, 97, 104, 94, 101, 104, 109, 106, 111, 105, 111, 111, 104, 94, 97, 128, 103, 113, 108, 114, 103, 103, 105, 97, 99, 108, 98, 107, 99, 95, 82, 104, 94, 73, 91, 109, 120, 146, 154, 155, 140, 124, 136, 142, 117, 118, 112, 89, 79, 92, 83, 88, 81, 80, 79, 80, 83, 77, 67, 50, 29, 20, 22, 53, 24, 31, 36, 31, 55, 49, 31, 13, 7, 0, 5, 7, 12, 15, 33, 40, 57, 82, 85, 86, 94, 93, 75, 93, 92, 102, 108, 115, 115, 112, 113, 122, 125, 109, 102, 97, 107, 110, 101, 117, 106, 111, 95, 94, 99, 128, 117, 112, 91, 104, 109, 115, 116, 104, 117, 100, 96, 92, 106, 113, 116, 108, 117, 110, 117, 109, 109, 118, 118, 119, 117, 123, 116, 117, 117, 117, 113, 123, 106, 119, 119, 122, 116, 118, 123, 120, 112, 112, 115, 119, 128, 124, 129, 132, 132, 131, 149, 133, 138, 142, 146, 140, 154, 155, 148, 142, 153, 145, 147, 152, 148, 151, 143, 142, 153, 153, 142, 149, 149, 153, 155, 154, 146, 149, 153, 137, 125, 120, 128, 127, 134, 133, 129, 124, 133, 126, 126, 133, 138, 132, 136, 124, 147, 140, 129, 137, 127, 127, 137, 135, 127, 101, 142, 119, 120, 120, 118, 120, 118, 110, 108, 97, 125, 127, 103, 92, 122, 94, 105, 101, 94, 82, 97, 106, 93, 116, 99, 84, 119, 111, 108, 101, 80, 89, 44, 86, 95, 47, 87, 97, 106, 108, 88, 71, 96, 89, 98, 103, 108, 106, 107, 111, 102, 106, 112, 109, 91, 117, 95, 108, 86, 81, 73, 152, 115, 102, 93, 109, 85, 98, 109, 115, 100, 107, 94, 79, 85, 122, 132, 154, 160, 160, 162, 157, 151, 146, 124, 118, 109, 80, 84, 81, 88, 86, 84, 89, 82, 76, 75, 79, 73, 62, 49, 37, 38, 64, 55, 46, 44, 32, 52, 74, 46, 14, 5, 11, 5, 12, 23, 36, 43, 50, 64, 71, 61, 72, 93, 81, 65, 85, 91, 101, 116, 124, 123, 115, 119, 116, 119, 103, 91, 93, 93, 99, 113, 114, 109, 102, 102, 105, 98, 117, 105, 110, 117, 111, 102, 110, 115, 97, 123, 107, 103, 99, 101, 107, 119, 100, 113, 112, 114, 117, 116, 113, 114, 110, 118, 110, 113, 108, 115, 117, 111, 117, 109, 121, 111, 122, 116, 121, 118, 114, 114, 118, 119, 118, 130, 127, 117, 129, 147, 127, 140, 143, 141, 126, 138, 148, 149, 143, 149, 147, 135, 114, 152, 160, 145, 151, 142, 137, 152, 153, 148, 148, 153, 149, 155, 143, 148, 148, 153, 157, 137, 139, 137, 129, 136, 131, 130, 124, 136, 122, 143, 134, 125, 137, 122, 115, 148, 150, 124, 132, 134, 119, 134, 133, 132, 121, 133, 118, 115, 120, 119, 113, 123, 116, 100, 98, 123, 117, 107, 99, 109, 101, 88, 81, 100, 66, 87, 113, 155, 122, 116, 115, 109, 101, 107, 105, 121, 22, 12, 73, 193, 75, 73, 90, 111, 86, 49, 99, 96, 78, 86, 107, 93, 112, 99, 108, 100, 101, 105, 107, 103, 114, 112, 109, 70, 79, 109, 147, 163, 107, 82, 100, 99, 92, 90, 127, 112, 109, 109, 95, 90, 124, 148, 161, 164, 163, 153, 127, 147, 172, 148, 117, 102, 95, 81, 60, 96, 119, 84, 87, 88, 74, 70, 68, 59, 56, 58, 46, 59, 51, 49, 50, 53, 58, 56, 75, 61, 31, 16, 15, 14, 24, 34, 41, 42, 59, 57, 60, 65, 76, 80, 71, 50, 70, 87, 95, 120, 119, 119, 119, 115, 107, 105, 99, 92, 93, 103, 107, 103, 107, 108, 110, 102, 105, 106, 114, 106, 111, 111, 114, 108, 106, 104, 113, 114, 111, 109, 116, 116, 109, 111, 103, 112, 116, 119, 120, 112, 105, 117, 117, 118, 110, 124, 109, 111, 108, 112, 108, 114, 111, 106, 108, 112, 108, 114, 116, 107, 132, 114, 123, 122, 127, 121, 134, 140, 130, 146, 139, 142, 139, 142, 128, 148, 145, 143, 148, 128, 111, 139, 152, 154, 144, 143, 149, 149, 152, 151, 158, 146, 139, 153, 147, 148, 140, 157, 157, 144, 138, 142, 129, 137, 137, 129, 127, 135, 126, 127, 136, 131, 138, 109, 95, 132, 154, 126, 129, 134, 126, 130, 132, 129, 130, 122, 130, 123, 124, 118, 117, 114, 123, 110, 112, 105, 118, 108, 109, 111, 102, 100, 79, 91, 106, 82, 83, 115, 144, 113, 115, 120, 105, 110, 114, 113, 0, 17, 50, 192, 127, 69, 101, 108, 21, 17, 114, 176, 88, 91, 96, 88, 111, 103, 101, 106, 111, 101, 90, 95, 121, 115, 98, 79, 71, 106, 140, 164, 118, 94, 108, 99, 90, 90, 107, 96, 85, 115, 96, 100, 132, 146, 159, 152, 149, 138, 113, 140, 169, 156, 105, 116, 98, 78, 60, 103, 96, 86, 83, 82, 79, 62, 65, 63, 60, 62, 47, 62, 49, 35, 59, 59, 43, 60, 78, 69, 38, 12, 20, 24, 32, 46, 39, 47, 56, 53, 59, 67, 75, 44, 92, 56, 68, 87, 100, 111, 113, 122, 113, 115, 113, 96, 95, 97, 99, 100, 107, 102, 107, 115, 108, 107, 112, 115, 108, 108, 111, 114, 109, 117, 113, 106, 105, 111, 113, 107, 111, 123, 115, 101, 108, 108, 122, 119, 122, 103, 113, 115, 116, 117, 117, 114, 109, 112, 91, 109, 114, 111, 113, 112, 120, 106, 116, 112, 116, 113, 124, 111, 123, 135, 134, 122, 135, 142, 130, 141, 135, 140, 143, 129, 127, 139, 142, 148, 149, 148, 145, 148, 150, 144, 144, 148, 148, 148, 146, 149, 148, 146, 148, 139, 148, 149, 154, 157, 154, 143, 131, 137, 132, 127, 132, 131, 138, 127, 129, 134, 127, 140, 133, 128, 108, 110, 131, 127, 133, 131, 131, 132, 135, 126, 126, 118, 131, 118, 127, 115, 118, 117, 114, 119, 116, 107, 117, 103, 117, 102, 108, 106, 52, 132, 98, 89, 112, 90, 103, 121, 116, 92, 107, 105, 107, 104, 33, 4, 43, 152, 117, 79, 109, 97, 33, 36, 75, 160, 78, 86, 101, 90, 96, 90, 106, 99, 111, 99, 102, 77, 112, 130, 107, 69, 74, 107, 124, 120, 126, 89, 105, 111, 103, 79, 68, 96, 80, 97, 99, 104, 141, 153, 160, 153, 146, 143, 113, 115, 138, 139, 93, 115, 98, 74, 62, 117, 96, 82, 98, 80, 79, 75, 79, 56, 77, 65, 61, 63, 22, 17, 65, 123, 83, 40, 64, 53, 45, 33, 24, 33, 43, 51, 52, 46, 39, 41, 84, 77, 75, 50, 59, 78, 65, 99, 104, 105, 121, 121, 112, 114, 104, 95, 103, 104, 99, 97, 111, 110, 106, 114, 104, 109, 109, 110, 114, 115, 107, 115, 104, 107, 119, 113, 104, 105, 112, 115, 118, 120, 121, 114, 107, 112, 115, 117, 114, 110, 115, 112, 112, 119, 122, 115, 110, 117, 108, 112, 103, 105, 126, 109, 108, 119, 122, 116, 118, 125, 126, 122, 129, 134, 130, 132, 131, 136, 134, 138, 134, 148, 136, 135, 143, 148, 150, 152, 145, 149, 143, 148, 153, 145, 144, 151, 152, 148, 139, 140, 149, 146, 144, 146, 154, 143, 157, 157, 153, 137, 131, 136, 137, 137, 127, 126, 127, 132, 127, 131, 131, 131, 127, 133, 136, 135, 130, 133, 135, 136, 127, 127, 130, 127, 124, 119, 121, 120, 130, 116, 119, 89, 116, 118, 117, 117, 114, 103, 102, 112, 109, 116, 58, 93, 119, 136, 124, 108, 109, 114, 115, 113, 111, 110, 98, 105, 92, 37, 53, 79, 86, 90, 101, 107, 90, 30, 45, 85, 76, 91, 88, 88, 91, 86, 101, 101, 101, 91, 95, 80, 103, 110, 118, 102, 88, 93, 105, 110, 103, 78, 89, 105, 95, 81, 84, 89, 75, 97, 95, 114, 126, 154, 169, 163, 153, 146, 132, 127, 126, 118, 93, 93, 99, 84, 53, 106, 119, 68, 107, 80, 82, 78, 73, 51, 93, 70, 75, 67, 13, 6, 55, 127, 97, 58, 63, 55, 42, 38, 38, 43, 52, 43, 47, 53, 44, 46, 78, 86, 67, 71, 95, 85, 86, 95, 98, 101, 103, 111, 111, 112, 103, 106, 100, 104, 102, 99, 105, 109, 112, 107, 117, 102, 106, 106, 114, 109, 108, 124, 121, 110, 121, 113, 110, 116, 112, 106, 116, 123, 117, 119, 120, 113, 125, 123, 112, 113, 118, 121, 115, 109, 122, 101, 108, 116, 115, 116, 99, 101, 131, 117, 108, 122, 124, 125, 118, 107, 104, 129, 127, 131, 134, 132, 125, 140, 131, 142, 143, 142, 141, 144, 146, 149, 146, 154, 144, 153, 150, 151, 149, 151, 149, 139, 153, 145, 147, 134, 152, 159, 142, 151, 146, 156, 139, 150, 144, 131, 127, 138, 138, 131, 125, 123, 136, 128, 131, 130, 131, 122, 125, 139, 128, 135, 131, 128, 131, 133, 127, 132, 131, 133, 118, 122, 121, 121, 126, 123, 114, 125, 124, 115, 116, 116, 113, 112, 107, 107, 124, 108, 103, 92, 89, 150, 97, 107, 116, 119, 123, 116, 111, 112, 112, 97, 103, 98, 87, 82, 100, 101, 76, 107, 95, 96, 83, 91, 113, 88, 89, 93, 86, 103, 97, 106, 95, 98, 105, 109, 107, 111, 109, 102, 112, 109, 98, 90, 106, 90, 100, 96, 87, 84, 88, 89, 88, 96, 102, 110, 112, 142, 160, 158, 160, 162, 145, 131, 124, 123, 111, 122, 93, 84, 60, 89, 105, 73, 75, 89, 79, 74, 75, 72, 75, 69, 81, 77, 41, 11, 46, 90, 67, 59, 68, 56, 43, 37, 66, 61, 59, 53, 49, 50, 57, 62, 82, 78, 71, 84, 94, 100, 91, 98, 98, 101, 104, 108, 116, 112, 104, 109, 107, 109, 106, 104, 115, 111, 109, 110, 114, 111, 103, 105, 118, 109, 114, 118, 109, 116, 117, 119, 108, 119, 121, 114, 124, 115, 125, 113, 115, 103, 129, 118, 104, 111, 115, 120, 119, 112, 115, 99, 117, 107, 113, 113, 99, 108, 115, 108, 109, 114, 118, 119, 113, 92, 104, 116, 114, 140, 139, 138, 131, 139, 135, 122, 172, 141, 141, 148, 145, 152, 146, 149, 150, 143, 153, 153, 151, 148, 154, 137, 154, 146, 146, 141, 149, 146, 142, 148, 144, 148, 143, 150, 146, 131, 138, 135, 137, 137, 137, 129, 129, 133, 128, 137, 129, 137, 127, 136, 144, 124, 138, 139, 129, 134, 126, 135, 131, 124, 125, 126, 114, 116, 138, 117, 117, 119, 129, 118, 107, 119, 113, 118, 107, 110, 104, 127, 124, 96, 68, 141, 119, 103, 118, 117, 113, 118, 101, 122, 109, 99, 107, 113, 96, 86, 107, 100, 96, 103, 86, 104, 98, 86, 89, 97, 89, 80, 100, 94, 103, 104, 68, 93, 127, 154, 95, 109, 103, 86, 120, 140, 109, 101, 102, 101, 128, 104, 93, 91, 83, 80, 93, 96, 85, 95, 120, 148, 160, 151, 149, 157, 147, 121, 120, 139, 130, 113, 69, 75, 128, 110, 93, 77, 58, 82, 76, 68, 72, 77, 72, 67, 61, 67, 94, 43, 48, 75, 69, 75, 67, 46, 38, 34, 60, 66, 65, 62, 59, 62, 65, 63, 74, 76, 83, 85, 102, 104, 96, 94, 95, 101, 100, 106, 118, 107, 103, 106, 105, 106, 110, 105, 117, 107, 124, 125, 110, 100, 108, 102, 107, 115, 122, 119, 122, 115, 114, 119, 120, 118, 123, 116, 124, 126, 120, 118, 106, 137, 114, 119, 122, 118, 108, 114, 109, 116, 106, 119, 114, 108, 108, 116, 118, 106, 110, 115, 106, 111, 107, 111, 113, 121, 99, 85, 119, 132, 141, 126, 136, 131, 131, 132, 147, 137, 148, 139, 151, 145, 155, 143, 145, 146, 150, 149, 153, 148, 157, 151, 148, 140, 149, 153, 149, 148, 145, 148, 148, 148, 146, 148, 146, 137, 127, 140, 138, 177, 140, 133, 129, 127, 124, 129, 131, 132, 127, 123, 139, 127, 131, 131, 130, 114, 125, 132, 131, 124, 126, 121, 125, 119, 116, 124, 126, 118, 128, 122, 114, 127, 109, 119, 108, 105, 107, 116, 116, 116, 91, 113, 107, 121, 120, 117, 121, 110, 113, 107, 104, 86, 123, 109, 110, 103, 99, 96, 104, 99, 97, 91, 96, 103, 89, 104, 83, 82, 87, 93, 97, 99, 66, 87, 127, 162, 104, 102, 99, 87, 109, 121, 96, 117, 93, 99, 121, 117, 105, 92, 88, 81, 85, 77, 84, 99, 122, 146, 159, 155, 154, 145, 130, 120, 105, 143, 130, 100, 48, 78, 146, 131, 90, 68, 75, 69, 67, 67, 60, 84, 72, 67, 38, 41, 98, 92, 58, 73, 75, 63, 54, 47, 48, 42, 51, 53, 78, 71, 71, 63, 46, 96, 69, 85, 86, 106, 99, 100, 96, 87, 80, 93, 92, 98, 110, 114, 105, 111, 107, 107, 112, 109, 116, 107, 121, 122, 106, 114, 101, 101, 107, 111, 113, 104, 117, 118, 121, 115, 120, 117, 121, 122, 118, 122, 113, 125, 109, 124, 115, 125, 118, 111, 115, 115, 105, 107, 116, 113, 114, 107, 100, 106, 111, 117, 116, 120, 108, 114, 120, 113, 124, 123, 115, 124, 119, 134, 136, 126, 138, 132, 142, 143, 143, 131, 146, 142, 148, 146, 143, 134, 152, 131, 151, 149, 149, 148, 151, 149, 155, 137, 156, 144, 153, 139, 146, 144, 157, 149, 151, 146, 157, 140, 124, 139, 137, 159, 137, 129, 128, 130, 133, 132, 125, 126, 136, 131, 129, 122, 130, 137, 131, 126, 131, 129, 124, 127, 127, 120, 128, 123, 122, 118, 116, 122, 122, 109, 117, 128, 116, 106, 107, 107, 111, 103, 101, 113, 119, 133, 112, 89, 115, 134, 116, 110, 112, 111, 105, 89, 109, 103, 100, 103, 114, 94, 100, 105, 91, 97, 109, 97, 95, 102, 79, 99, 100, 95, 101, 104, 77, 86, 112, 124, 107, 116, 114, 107, 107, 105, 101, 111, 109, 110, 108, 95, 111, 96, 108, 90, 90, 66, 80, 98, 118, 132, 139, 166, 163, 137, 132, 130, 137, 157, 124, 97, 60, 68, 119, 107, 84, 53, 93, 102, 65, 84, 60, 75, 65, 51, 39, 49, 68, 71, 64, 66, 82, 71, 56, 47, 54, 46, 53, 61, 73, 75, 81, 76, 58, 73, 80, 97, 107, 102, 91, 88, 91, 83, 78, 87, 90, 93, 103, 112, 107, 111, 117, 109, 116, 120, 110, 116, 110, 113, 111, 108, 106, 84, 114, 109, 114, 119, 123, 111, 120, 114, 126, 117, 121, 110, 124, 143, 111, 114, 125, 124, 121, 114, 119, 117, 110, 109, 112, 107, 110, 119, 108, 94, 106, 106, 117, 113, 107, 115, 117, 115, 114, 125, 123, 125, 128, 138, 124, 137, 130, 128, 136, 127, 136, 151, 142, 137, 151, 144, 148, 138, 146, 149, 143, 146, 149, 146, 143, 148, 148, 144, 141, 142, 148, 141, 146, 140, 155, 148, 151, 139, 150, 146, 150, 137, 133, 137, 131, 147, 141, 135, 134, 131, 132, 131, 136, 129, 140, 132, 139, 116, 141, 131, 133, 128, 130, 129, 129, 127, 129, 127, 124, 121, 117, 125, 115, 124, 128, 114, 119, 120, 123, 121, 112, 113, 113, 116, 104, 92, 114, 137, 118, 102, 103, 116, 101, 110, 99, 128, 103, 100, 102, 104, 103, 107, 94, 93, 102, 95, 94, 91, 101, 92, 106, 100, 97, 90, 103, 104, 100, 106, 98, 94, 104, 114, 92, 113, 109, 106, 111, 115, 106, 110, 110, 121, 114, 97, 90, 95, 117, 93, 81, 89, 87, 93, 106, 105, 104, 145, 158, 136, 132, 145, 143, 161, 147, 108, 107, 91, 107, 86, 63, 35, 72, 85, 71, 88, 68, 71, 66, 61, 52, 75, 79, 71, 61, 66, 68, 65, 57, 53, 54, 53, 52, 72, 78, 83, 78, 72, 75, 77, 101, 104, 108, 106, 99, 93, 95, 88, 74, 80, 79, 88, 96, 113, 109, 116, 114, 108, 116, 111, 113, 117, 117, 107, 110, 109, 108, 107, 109, 109, 116, 128, 119, 117, 120, 118, 119, 124, 117, 110, 112, 139, 123, 122, 125, 120, 133, 115, 119, 125, 117, 112, 112, 109, 110, 114, 116, 109, 108, 118, 114, 116, 117, 122, 121, 124, 111, 126, 129, 127, 126, 137, 134, 137, 132, 135, 145, 110, 122, 166, 150, 140, 146, 142, 139, 152, 143, 149, 152, 156, 147, 153, 143, 155, 148, 156, 146, 142, 144, 148, 142, 146, 145, 142, 153, 146, 134, 142, 149, 138, 135, 144, 131, 155, 133, 129, 131, 126, 137, 131, 127, 133, 128, 126, 128, 127, 118, 130, 138, 134, 137, 129, 123, 129, 126, 124, 127, 119, 124, 127, 127, 122, 136, 115, 125, 119, 120, 115, 109, 117, 110, 113, 108, 96, 127, 120, 103, 114, 112, 118, 114, 105, 95, 124, 89, 107, 108, 102, 97, 98, 90, 86, 103, 92, 88, 99, 103, 98, 101, 107, 98, 96, 104, 98, 102, 107, 106, 102, 107, 116, 104, 103, 108, 115, 117, 106, 108, 114, 118, 108, 112, 105, 85, 95, 121, 109, 97, 89, 98, 90, 108, 104, 95, 103, 135, 124, 136, 153, 152, 160, 168, 152, 137, 123, 105, 97, 75, 56, 52, 65, 57, 80, 75, 74, 61, 69, 66, 52, 84, 62, 53, 66, 66, 66, 59, 64, 60, 60, 59, 75, 76, 67, 74, 71, 83, 90, 114, 118, 121, 108, 110, 100, 87, 84, 78, 76, 75, 88, 100, 115, 102, 113, 112, 113, 118, 117, 119, 116, 122, 115, 115, 109, 111, 121, 111, 113, 120, 122, 122, 125, 116, 126, 118, 125, 124, 126, 110, 105, 124, 148, 124, 118, 127, 117, 119, 117, 121, 119, 115, 117, 109, 106, 112, 119, 104, 125, 133, 119, 120, 116, 119, 127, 121, 127, 130, 131, 125, 129, 141, 139, 136, 114, 125, 129, 123, 141, 140, 135, 141, 138, 142, 145, 136, 146, 153, 150, 146, 144, 150, 155, 146, 148, 148, 146, 144, 142, 156, 146, 146, 140, 149, 146, 149, 149, 132, 137, 129, 148, 190, 142, 129, 127, 143, 126, 131, 132, 131, 133, 113, 117, 129, 121, 114, 123, 135, 129, 127, 133, 127, 118, 126, 130, 125, 124, 126, 120, 130, 115, 124, 127, 132, 119, 118, 108, 140, 108, 111, 122, 119, 106, 115, 94, 117, 109, 106, 108, 116, 87, 103, 128, 83, 103, 118, 90, 99, 96, 103, 96, 98, 90, 94, 93, 91, 99, 103, 101, 100, 90, 89, 103, 102, 117, 100, 114, 112, 114, 120, 98, 109, 117, 109, 110, 113, 117, 111, 106, 103, 107, 90, 93, 91, 120, 105, 99, 100, 100, 110, 110, 89, 93, 110, 119, 124, 155, 156, 158, 162, 171, 159, 127, 121, 111, 86, 82, 61, 63, 68, 66, 70, 70, 69, 61, 66, 61, 78, 46, 31, 53, 66, 66, 67, 65, 56, 54, 70, 77, 74, 66, 71, 84, 100, 108, 102, 112, 118, 122, 113, 93, 80, 80, 75, 65, 66, 81, 103, 111, 116, 118, 118, 120, 107, 116, 115, 116, 111, 97, 117, 120, 114, 114, 116, 122, 121, 111, 120, 120, 113, 119, 120, 121, 127, 123, 119, 104, 131, 134, 121, 131, 123, 118, 124, 118, 126, 118, 111, 109, 107, 114, 98, 115, 105, 127, 131, 116, 129, 120, 116, 123, 121, 127, 120, 93, 106, 120, 138, 137, 124, 143, 128, 132, 138, 137, 131, 145, 135, 139, 140, 141, 154, 148, 141, 156, 147, 147, 148, 147, 148, 151, 155, 146, 145, 149, 141, 146, 146, 144, 137, 151, 148, 146, 146, 138, 141, 131, 146, 140, 129, 126, 135, 133, 130, 110, 131, 122, 131, 126, 126, 126, 126, 124, 125, 127, 127, 132, 123, 129, 124, 127, 124, 130, 126, 119, 132, 124, 127, 117, 114, 122, 114, 86, 128, 115, 111, 109, 107, 113, 116, 104, 112, 112, 101, 104, 107, 92, 110, 109, 87, 92, 124, 89, 98, 93, 96, 94, 91, 94, 97, 103, 106, 92, 94, 102, 98, 95, 104, 106, 106, 110, 100, 108, 102, 107, 122, 106, 110, 109, 111, 109, 107, 104, 113, 111, 109, 102, 95, 99, 98, 96, 105, 105, 103, 102, 110, 114, 80, 97, 109, 100, 103, 146, 152, 160, 167, 167, 176, 142, 124, 109, 95, 84, 67, 81, 77, 62, 73, 80, 77, 63, 68, 62, 69, 52, 36, 48, 57, 69, 74, 73, 50, 55, 87, 85, 84, 73, 74, 85, 109, 109, 112, 115, 120, 121, 100, 88, 76, 78, 70, 66, 60, 87, 97, 111, 121, 114, 99, 104, 121, 115, 125, 114, 107, 95, 122, 139, 121, 126, 120, 114, 110, 119, 115, 125, 120, 117, 117, 122, 132, 128, 128, 122, 126, 127, 124, 121, 123, 124, 123, 120, 127, 122, 122, 109, 112, 104, 114, 118, 104, 123, 108, 109, 120, 122, 113, 127, 116, 111, 125, 122, 107, 128, 133, 133, 119, 140, 137, 143, 139, 128, 140, 137, 130, 146, 142, 146, 146, 149, 136, 148, 134, 140, 146, 141, 151, 151, 151, 149, 146, 144, 148, 141, 138, 140, 147, 149, 140, 143, 155, 137, 131, 127, 137, 131, 125, 136, 123, 146, 129, 124, 129, 129, 131, 127, 126, 133, 129, 126, 129, 122, 118, 137, 127, 124, 121, 134, 122, 118, 126, 121, 126, 121, 114, 126, 121, 124, 118, 119, 121, 121, 109, 113, 118, 114, 114, 110, 111, 121, 102, 87, 113, 95, 115, 112, 102, 112, 103, 90, 102, 94, 95, 86, 88, 109, 98, 108, 102, 102, 104, 79, 117, 108, 97, 103, 105, 117, 106, 117, 112, 111, 117, 119, 115, 109, 109, 105, 90, 104, 107, 111, 113, 107, 90, 95, 94, 110, 101, 100, 100, 87, 107, 113, 97, 97, 87, 42, 69, 116, 133, 147, 161, 171, 164, 148, 130, 108, 94, 88, 80, 82, 79, 69, 71, 75, 74, 67, 62, 60, 69, 56, 57, 50, 55, 57, 78, 80, 47, 42, 84, 89, 90, 79, 70, 89, 105, 104, 114, 118, 119, 115, 107, 94, 79, 83, 78, 65, 66, 75, 95, 117, 116, 113, 111, 104, 117, 121, 122, 114, 114, 101, 122, 116, 112, 114, 107, 109, 99, 114, 107, 108, 127, 117, 118, 116, 134, 128, 129, 127, 126, 127, 117, 122, 123, 128, 127, 121, 119, 117, 121, 121, 112, 107, 112, 123, 122, 121, 121, 108, 115, 121, 135, 145, 122, 122, 119, 128, 123, 134, 136, 132, 138, 134, 137, 135, 147, 139, 139, 123, 124, 137, 147, 141, 138, 147, 140, 155, 137, 136, 148, 153, 153, 145, 148, 153, 149, 146, 144, 148, 146, 138, 140, 146, 140, 148, 153, 140, 140, 122, 135, 133, 126, 123, 132, 129, 118, 127, 127, 131, 129, 127, 130, 135, 133, 131, 134, 131, 131, 133, 124, 136, 126, 129, 122, 124, 127, 129, 128, 116, 107, 125, 119, 118, 119, 111, 96, 110, 123, 109, 114, 116, 117, 116, 109, 110, 107, 93, 109, 92, 101, 96, 102, 105, 100, 77, 120, 98, 83, 76, 90, 96, 106, 103, 100, 91, 90, 103, 99, 98, 108, 115, 115, 106, 102, 110, 112, 106, 106, 109, 109, 114, 112, 104, 105, 111, 108, 104, 107, 102, 104, 81, 91, 102, 102, 102, 102, 123, 103, 98, 107, 111, 96, 68, 71, 92, 117, 144, 157, 160, 154, 131, 124, 112, 102, 85, 80, 86, 82, 75, 64, 81, 64, 67, 64, 66, 71, 79, 70, 64, 67, 63, 95, 88, 75, 69, 80, 92, 90, 88, 81, 92, 103, 102, 103, 105, 119, 115, 111, 95, 90, 86, 77, 76, 74, 85, 94, 123, 128, 121, 115, 108, 113, 118, 117, 120, 125, 118, 124, 119, 114, 117, 114, 105, 85, 93, 112, 115, 120, 116, 123, 115, 125, 122, 130, 127, 120, 120, 122, 118, 131, 130, 129, 124, 115, 126, 117, 114, 120, 112, 88, 119, 112, 117, 119, 112, 114, 114, 123, 131, 122, 114, 123, 133, 129, 135, 140, 131, 138, 130, 147, 136, 141, 142, 137, 134, 147, 136, 142, 148, 144, 139, 138, 149, 142, 147, 154, 147, 151, 149, 153, 143, 151, 144, 142, 142, 135, 146, 142, 137, 151, 144, 148, 133, 131, 122, 133, 121, 143, 124, 125, 131, 116, 143, 126, 129, 127, 140, 129, 131, 129, 130, 127, 133, 131, 134, 136, 124, 116, 131, 111, 119, 122, 132, 129, 123, 125, 119, 108, 120, 109, 112, 110, 118, 113, 103, 114, 113, 113, 111, 112, 114, 94, 108, 110, 99, 109, 98, 102, 103, 90, 87, 89, 100, 92, 84, 100, 101, 98, 79, 129, 96, 97, 98, 110, 108, 104, 105, 100, 117, 112, 107, 122, 115, 112, 107, 107, 108, 103, 113, 112, 116, 117, 105, 102, 106, 107, 94, 104, 115, 93, 102, 103, 101, 109, 104, 113, 123, 113, 91, 80, 84, 98, 126, 149, 146, 137, 134, 146, 100, 87, 86, 68, 90, 84, 82, 73, 69, 75, 80, 73, 74, 77, 86, 77, 64, 61, 58, 86, 87, 88, 89, 86, 99, 93, 96, 94, 96, 107, 113, 116, 117, 115, 113, 105, 89, 80, 87, 83, 69, 69, 94, 104, 113, 123, 119, 117, 117, 118, 124, 125, 118, 125, 124, 124, 123, 112, 120, 121, 115, 99, 107, 106, 120, 128, 117, 119, 118, 124, 118, 119, 129, 122, 125, 124, 121, 123, 138, 124, 127, 118, 123, 124, 125, 118, 119, 108, 120, 121, 112, 121, 120, 117, 109, 125, 120, 121, 122, 122, 122, 130, 132, 134, 137, 140, 140, 141, 135, 137, 139, 131, 142, 138, 141, 142, 141, 140, 142, 140, 145, 146, 143, 143, 146, 146, 138, 136, 147, 151, 149, 138, 157, 138, 140, 146, 133, 149, 140, 140, 135, 131, 126, 126, 125, 126, 127, 127, 131, 108, 126, 104, 138, 120, 127, 124, 120, 127, 116, 135, 131, 133, 127, 133, 128, 121, 126, 111, 110, 126, 128, 122, 123, 115, 109, 119, 115, 111, 118, 113, 108, 107, 104, 103, 111, 112, 111, 108, 107, 94, 105, 109, 107, 90, 103, 92, 119, 100, 105, 89, 97, 97, 99, 101, 100, 105, 77, 109, 98, 85, 95, 107, 110, 106, 114, 108, 107, 109, 105, 124, 114, 117, 111, 103, 92, 100, 97, 104, 115, 108, 83, 86, 105, 101, 84, 97, 118, 85, 74, 108, 99, 104, 113, 115, 122, 109, 104, 100, 84, 93, 109, 127, 136, 125, 121, 129, 100, 84, 87, 80, 91, 87, 81, 76, 72, 77, 78, 75, 86, 83, 76, 73, 79, 82, 74, 87, 91, 94, 89, 93, 92, 88, 96, 93, 89, 104, 121, 119, 115, 111, 107, 91, 84, 76, 84, 74, 61, 84, 110, 111, 113, 115, 113, 118, 117, 115, 125, 123, 122, 127, 115, 125, 120, 119, 117, 125, 113, 112, 118, 115, 115, 120, 121, 121, 125, 125, 117, 121, 122, 119, 125, 122, 118, 129, 132, 124, 124, 127, 117, 125, 121, 122, 124, 118, 128, 116, 112, 110, 119, 123, 105, 108, 126, 125, 125, 139, 130, 127, 132, 128, 126, 147, 138, 128, 139, 129, 131, 133, 144, 130, 125, 140, 135, 128, 141, 146, 141, 150, 146, 142, 148, 144, 142, 117, 139, 155, 141, 142, 147, 140, 132, 151, 155, 147, 134, 149, 135, 127, 148, 137, 118, 127, 131, 124, 117, 113, 120, 118, 122, 118, 117, 124, 115, 120, 111, 130, 129, 136, 127, 125, 133, 131, 115, 118, 124, 127, 128, 124, 119, 116, 116, 113, 117, 99, 112, 99, 97, 106, 107, 109, 109, 111, 117, 112, 103, 112, 109, 105, 108, 105, 98, 89, 104, 100, 96, 108, 95, 99, 100, 95, 104, 107, 100, 105, 91, 103, 95, 100, 106, 109, 100, 106, 115, 115, 112, 118, 119, 112, 119, 73, 63, 154, 132, 100, 112, 106, 94, 98, 72, 49, 117, 96, 109, 99, 93, 95, 101, 114, 118, 108, 125, 116, 104, 108, 90, 91, 90, 104, 126, 120, 123, 106, 95, 73, 73, 83, 97, 104, 84, 76, 76, 84, 93, 87, 81, 78, 77, 77, 88, 90, 86, 86, 81, 81, 108, 105, 96, 82, 92, 85, 99, 117, 118, 114, 115, 110, 91, 78, 68, 74, 82, 83, 88, 103, 118, 117, 117, 112, 117, 123, 121, 123, 123, 122, 125, 120, 124, 124, 126, 129, 115, 113, 113, 118, 119, 113, 116, 124, 123, 123, 127, 123, 117, 125, 118, 115, 131, 128, 127, 128, 124, 122, 123, 122, 120, 124, 119, 116, 118, 119, 128, 125, 118, 97, 94, 121, 119, 126, 139, 147, 122, 120, 135, 134, 128, 140, 121, 141, 145, 136, 130, 139, 137, 136, 140, 133, 136, 135, 146, 145, 144, 138, 140, 154, 145, 154, 148, 141, 142, 140, 151, 148, 148, 136, 140, 146, 135, 148, 146, 144, 151, 142, 131, 124, 126, 129, 124, 127, 129, 122, 122, 118, 120, 124, 117, 111, 104, 120, 87, 113, 111, 120, 124, 119, 150, 124, 131, 129, 126, 129, 117, 121, 126, 120, 124, 120, 123, 103, 125, 126, 112, 103, 97, 106, 107, 111, 108, 108, 114, 111, 106, 113, 97, 98, 119, 103, 110, 93, 101, 96, 70, 100, 110, 87, 93, 88, 95, 101, 99, 104, 99, 99, 102, 104, 103, 109, 103, 104, 112, 111, 116, 123, 106, 121, 114, 54, 49, 153, 148, 100, 108, 116, 113, 105, 40, 29, 120, 100, 102, 114, 106, 110, 108, 109, 117, 114, 116, 107, 99, 106, 93, 77, 73, 118, 153, 120, 131, 104, 89, 89, 81, 83, 86, 93, 88, 86, 81, 84, 92, 87, 84, 67, 75, 83, 87, 91, 77, 76, 77, 89, 108, 98, 98, 86, 77, 54, 98, 127, 113, 107, 106, 92, 73, 70, 59, 56, 74, 83, 99, 108, 113, 118, 109, 115, 118, 117, 116, 117, 121, 126, 113, 118, 135, 127, 125, 126, 121, 119, 120, 119, 119, 110, 120, 127, 130, 122, 121, 126, 127, 125, 120, 108, 130, 123, 121, 125, 128, 117, 123, 119, 122, 124, 118, 123, 116, 122, 121, 122, 119, 117, 119, 119, 120, 127, 132, 140, 143, 140, 141, 133, 135, 139, 126, 137, 148, 136, 130, 136, 141, 124, 137, 134, 142, 147, 141, 139, 144, 144, 153, 139, 134, 139, 155, 138, 152, 146, 149, 148, 142, 151, 150, 148, 140, 138, 146, 137, 151, 140, 140, 124, 131, 129, 126, 129, 131, 122, 117, 122, 122, 118, 115, 117, 109, 110, 109, 111, 113, 120, 125, 102, 147, 124, 131, 116, 130, 127, 131, 122, 129, 118, 117, 104, 110, 126, 114, 111, 113, 105, 106, 99, 112, 113, 109, 110, 114, 107, 105, 118, 105, 93, 111, 106, 90, 112, 97, 103, 74, 95, 103, 97, 91, 89, 106, 101, 96, 93, 100, 98, 105, 103, 110, 111, 107, 117, 120, 102, 119, 117, 104, 140, 122, 88, 52, 104, 108, 102, 115, 116, 113, 113, 69, 55, 102, 95, 111, 99, 98, 102, 114, 92, 127, 119, 113, 90, 90, 100, 74, 69, 53, 131, 137, 130, 123, 102, 95, 93, 87, 85, 89, 82, 92, 97, 88, 87, 76, 84, 89, 69, 70, 105, 91, 81, 89, 84, 84, 79, 90, 95, 112, 115, 99, 84, 97, 127, 114, 107, 106, 80, 66, 66, 56, 47, 66, 83, 94, 120, 118, 110, 119, 123, 110, 127, 125, 120, 112, 126, 128, 118, 130, 115, 124, 128, 119, 121, 119, 114, 122, 112, 117, 120, 120, 123, 121, 124, 127, 125, 126, 122, 129, 117, 115, 124, 129, 120, 120, 123, 130, 118, 122, 113, 123, 121, 125, 130, 126, 123, 125, 116, 123, 127, 129, 134, 133, 126, 159, 149, 138, 126, 142, 132, 128, 146, 135, 130, 132, 109, 101, 137, 132, 127, 133, 146, 140, 140, 142, 148, 141, 141, 145, 140, 142, 138, 148, 144, 141, 146, 155, 146, 144, 142, 140, 142, 142, 142, 133, 131, 124, 133, 126, 133, 126, 123, 120, 129, 107, 105, 118, 115, 113, 115, 112, 112, 118, 115, 113, 128, 131, 133, 124, 124, 126, 124, 128, 122, 119, 118, 117, 116, 109, 123, 117, 108, 108, 112, 104, 109, 111, 113, 112, 105, 111, 109, 109, 104, 104, 107, 100, 105, 82, 113, 90, 113, 97, 97, 98, 92, 78, 121, 90, 103, 109, 107, 89, 106, 103, 113, 111, 107, 112, 119, 121, 114, 118, 122, 110, 121, 113, 117, 96, 99, 77, 114, 114, 121, 118, 120, 103, 87, 122, 98, 110, 105, 99, 106, 115, 117, 115, 122, 104, 79, 114, 84, 64, 67, 71, 106, 116, 137, 132, 119, 104, 96, 85, 77, 77, 96, 100, 94, 94, 90, 93, 91, 86, 47, 58, 143, 110, 80, 86, 84, 93, 89, 76, 89, 108, 117, 122, 101, 100, 120, 120, 110, 91, 71, 62, 52, 57, 54, 62, 83, 103, 118, 115, 113, 117, 120, 113, 127, 123, 116, 98, 123, 127, 126, 122, 115, 122, 137, 121, 115, 120, 124, 119, 119, 120, 125, 109, 128, 114, 114, 121, 118, 130, 128, 126, 125, 126, 128, 127, 119, 132, 119, 124, 121, 113, 122, 120, 124, 127, 135, 127, 127, 121, 120, 123, 129, 125, 127, 122, 134, 133, 140, 146, 131, 133, 131, 127, 129, 129, 137, 131, 112, 105, 132, 123, 130, 142, 146, 150, 136, 137, 143, 147, 144, 137, 134, 146, 144, 148, 152, 142, 155, 144, 148, 138, 140, 129, 144, 149, 144, 137, 131, 131, 118, 131, 126, 117, 115, 120, 111, 107, 115, 115, 113, 117, 117, 113, 103, 127, 120, 112, 126, 119, 129, 126, 122, 126, 124, 124, 122, 124, 125, 122, 111, 109, 115, 114, 102, 94, 97, 109, 111, 107, 106, 112, 107, 114, 103, 96, 109, 110, 95, 111, 103, 97, 107, 85, 92, 114, 95, 100, 77, 105, 95, 111, 115, 107, 100, 104, 105, 105, 114, 113, 111, 119, 126, 118, 101, 108, 118, 116, 122, 119, 116, 119, 107, 106, 108, 112, 116, 113, 109, 105, 87, 92, 97, 98, 105, 111, 101, 108, 104, 122, 112, 104, 87, 97, 73, 54, 66, 92, 113, 115, 131, 132, 115, 103, 102, 92, 70, 73, 86, 78, 62, 114, 148, 106, 89, 87, 60, 53, 112, 98, 77, 92, 98, 95, 100, 93, 86, 86, 104, 119, 113, 107, 110, 108, 91, 80, 68, 54, 40, 58, 60, 76, 82, 97, 76, 140, 104, 117, 118, 104, 130, 147, 117, 122, 113, 125, 131, 125, 115, 118, 136, 126, 120, 122, 123, 130, 127, 123, 124, 122, 120, 103, 116, 117, 121, 120, 130, 124, 122, 126, 130, 127, 132, 128, 122, 130, 130, 119, 125, 125, 130, 130, 127, 127, 112, 129, 109, 118, 126, 135, 132, 121, 122, 138, 128, 137, 127, 128, 124, 113, 139, 127, 129, 135, 133, 125, 132, 137, 126, 143, 142, 152, 139, 143, 146, 144, 137, 126, 144, 151, 144, 135, 148, 144, 153, 144, 144, 142, 148, 127, 142, 142, 146, 131, 117, 133, 133, 124, 120, 109, 107, 124, 119, 98, 120, 120, 122, 111, 121, 113, 115, 124, 123, 114, 126, 113, 141, 126, 120, 126, 124, 122, 118, 133, 124, 121, 112, 107, 107, 107, 91, 83, 91, 93, 104, 111, 92, 111, 108, 102, 104, 92, 102, 89, 98, 97, 108, 88, 96, 98, 97, 88, 101, 99, 96, 99, 97, 106, 105, 96, 106, 106, 120, 111, 112, 105, 114, 125, 114, 116, 107, 109, 112, 114, 122, 120, 105, 121, 104, 105, 112, 108, 107, 119, 108, 102, 107, 96, 93, 95, 98, 106, 104, 90, 97, 106, 114, 112, 104, 102, 76, 66, 76, 92, 107, 119, 132, 121, 104, 99, 105, 100, 83, 83, 84, 55, 62, 114, 126, 100, 83, 79, 85, 79, 88, 68, 76, 92, 104, 95, 98, 101, 92, 88, 102, 110, 110, 126, 115, 108, 101, 71, 55, 50, 53, 56, 67, 80, 85, 101, 74, 127, 82, 110, 122, 93, 128, 140, 125, 124, 121, 118, 130, 122, 137, 123, 129, 119, 116, 114, 131, 127, 121, 123, 120, 119, 121, 95, 116, 114, 125, 118, 124, 118, 118, 123, 118, 125, 122, 121, 124, 126, 133, 122, 126, 126, 119, 126, 120, 127, 123, 124, 129, 124, 133, 127, 133, 128, 119, 134, 134, 134, 127, 123, 122, 117, 127, 129, 132, 130, 125, 129, 135, 140, 137, 147, 146, 142, 147, 147, 146, 148, 142, 145, 142, 142, 146, 153, 140, 144, 155, 146, 140, 138, 148, 135, 149, 133, 146, 133, 122, 126, 127, 126, 118, 124, 113, 124, 117, 126, 122, 117, 115, 111, 127, 122, 120, 103, 136, 111, 113, 117, 124, 123, 125, 122, 127, 124, 121, 117, 114, 116, 115, 117, 113, 108, 100, 73, 93, 95, 104, 104, 98, 97, 100, 102, 101, 96, 101, 99, 103, 95, 105, 93, 91, 96, 96, 97, 97, 101, 89, 116, 99, 105, 112, 99, 99, 104, 116, 109, 107, 109, 114, 127, 106, 114, 126, 107, 113, 109, 113, 125, 93, 103, 110, 111, 109, 110, 120, 114, 106, 113, 109, 103, 83, 88, 98, 97, 104, 96, 90, 108, 115, 105, 99, 93, 89, 81, 80, 86, 90, 103, 119, 109, 84, 84, 108, 116, 120, 112, 93, 71, 61, 83, 93, 80, 78, 88, 82, 75, 95, 93, 83, 92, 87, 97, 95, 105, 106, 89, 108, 122, 124, 107, 103, 107, 93, 39, 36, 44, 48, 46, 65, 76, 84, 108, 125, 109, 105, 108, 130, 120, 122, 123, 116, 129, 122, 128, 128, 127, 128, 123, 123, 121, 123, 120, 127, 125, 124, 128, 116, 119, 119, 106, 111, 114, 116, 104, 121, 135, 132, 122, 129, 132, 123, 121, 121, 120, 128, 122, 121, 127, 129, 131, 133, 131, 126, 129, 123, 123, 126, 131, 133, 131, 130, 141, 137, 138, 138, 136, 130, 127, 126, 136, 143, 136, 132, 137, 137, 135, 129, 136, 139, 148, 148, 139, 144, 142, 134, 131, 155, 135, 148, 142, 144, 149, 148, 142, 142, 146, 140, 131, 144, 142, 146, 129, 127, 133, 126, 127, 129, 124, 126, 117, 107, 144, 126, 120, 120, 122, 126, 127, 123, 96, 136, 146, 105, 121, 123, 119, 127, 129, 122, 124, 122, 121, 115, 102, 116, 101, 106, 112, 96, 87, 88, 103, 107, 106, 98, 92, 96, 105, 104, 97, 96, 101, 102, 101, 102, 114, 92, 103, 79, 88, 95, 98, 99, 115, 110, 95, 112, 101, 109, 103, 112, 109, 111, 117, 113, 129, 108, 128, 113, 102, 114, 118, 97, 117, 118, 116, 119, 106, 101, 89, 106, 103, 87, 112, 110, 106, 91, 78, 90, 80, 99, 96, 84, 109, 107, 97, 93, 102, 93, 90, 94, 97, 86, 93, 88, 98, 83, 86, 95, 108, 128, 126, 106, 99, 90, 90, 99, 88, 81, 74, 69, 83, 91, 88, 84, 88, 92, 96, 87, 102, 112, 109, 103, 123, 127, 110, 105, 94, 91, 69, 51, 43, 50, 54, 60, 76, 82, 103, 121, 118, 128, 113, 115, 128, 123, 122, 123, 128, 120, 132, 127, 127, 128, 126, 127, 128, 121, 119, 122, 126, 126, 114, 115, 115, 127, 122, 112, 120, 109, 119, 111, 129, 146, 130, 131, 132, 129, 124, 120, 122, 127, 110, 126, 147, 130, 125, 129, 131, 131, 121, 131, 127, 127, 128, 124, 132, 133, 136, 138, 135, 133, 136, 134, 136, 142, 142, 143, 129, 142, 138, 148, 130, 141, 134, 148, 142, 142, 138, 161, 142, 133, 140, 140, 135, 148, 142, 142, 142, 144, 144, 144, 142, 140, 137, 131, 146, 135, 111, 127, 127, 124, 133, 129, 131, 126, 129, 122, 131, 124, 135, 128, 115, 129, 131, 126, 82, 101, 159, 125, 115, 114, 123, 116, 112, 120, 117, 112, 122, 118, 104, 97, 93, 100, 115, 101, 99, 102, 98, 108, 109, 105, 93, 108, 107, 105, 107, 84, 101, 98, 94, 87, 104, 98, 97, 93, 104, 99, 88, 110, 112, 92, 99, 107, 90, 114, 122, 106, 109, 106, 123, 121, 150, 106, 118, 117, 116, 109, 107, 109, 110, 91, 122, 109, 102, 103, 100, 94, 97, 97, 103, 106, 107, 97, 89, 86, 87, 89, 94, 95, 100, 91, 93, 84, 97, 103, 83, 93, 96, 77, 94, 92, 74, 79, 93, 96, 98, 110, 103, 99, 123, 104, 96, 105, 93, 93, 85, 78, 86, 90, 82, 88, 88, 100, 99, 98, 91, 101, 113, 108, 121, 123, 117, 108, 97, 100, 77, 57, 53, 54, 51, 66, 74, 87, 102, 108, 105, 129, 120, 110, 130, 138, 123, 127, 126, 121, 121, 123, 125, 127, 130, 132, 130, 125, 125, 125, 124, 126, 125, 125, 113, 131, 117, 108, 118, 102, 117, 121, 119, 129, 107, 131, 139, 124, 134, 122, 129, 136, 126, 130, 128, 124, 125, 128, 128, 137, 102, 144, 126, 122, 130, 128, 134, 133, 135, 135, 134, 138, 135, 135, 134, 118, 138, 145, 130, 143, 120, 150, 133, 144, 139, 137, 147, 118, 141, 174, 135, 138, 140, 140, 144, 156, 148, 153, 138, 140, 146, 142, 138, 148, 148, 137, 146, 142, 133, 131, 133, 127, 129, 129, 127, 127, 126, 138, 131, 131, 127, 129, 133, 133, 136, 127, 108, 100, 128, 121, 108, 128, 126, 125, 115, 115, 111, 115, 116, 107, 129, 106, 107, 108, 95, 91, 97, 104, 109, 99, 114, 103, 105, 111, 114, 106, 106, 101, 103, 102, 97, 80, 86, 102, 89, 98, 94, 101, 96, 104, 96, 109, 99, 112, 104, 105, 108, 111, 112, 110, 110, 118, 128, 125, 112, 116, 118, 110, 102, 114, 116, 102, 107, 107, 106, 107, 95, 102, 105, 109, 105, 101, 105, 101, 95, 85, 88, 84, 99, 83, 93, 93, 84, 84, 95, 98, 88, 97, 90, 88, 98, 98, 98, 108, 97, 95, 95, 72, 67, 80, 134, 133, 115, 104, 94, 94, 86, 85, 92, 94, 88, 92, 95, 103, 93, 86, 88, 100, 93, 101, 125, 122, 117, 113, 102, 92, 70, 56, 52, 53, 57, 69, 71, 81, 93, 110, 102, 117, 110, 115, 125, 132, 126, 129, 125, 127, 115, 126, 120, 129, 135, 125, 134, 128, 125, 128, 123, 132, 127, 140, 165, 127, 105, 94, 115, 123, 118, 118, 122, 128, 124, 125, 129, 125, 137, 130, 118, 121, 125, 134, 124, 125, 121, 119, 134, 134, 132, 132, 120, 124, 131, 127, 131, 131, 133, 126, 129, 143, 139, 140, 134, 131, 137, 146, 137, 142, 121, 144, 147, 134, 146, 145, 152, 113, 135, 153, 146, 144, 146, 138, 132, 143, 146, 148, 142, 146, 144, 149, 151, 138, 142, 138, 149, 149);
constant memory:MEM_array:=(150, 144, 155, 157, 105, 164, 173, 173, 171, 173, 177, 181, 178, 183, 178, 180, 184, 186, 190, 183, 185, 185, 184, 188, 188, 185, 183, 190, 187, 187, 188, 186, 190, 189, 190, 190, 190, 192, 193, 193, 193, 192, 191, 194, 197, 195, 198, 196, 194, 193, 193, 196, 194, 199, 198, 200, 198, 198, 195, 195, 196, 200, 200, 198, 199, 199, 200, 197, 198, 199, 203, 198, 202, 200, 200, 200, 200, 201, 201, 200, 202, 199, 200, 201, 203, 199, 204, 201, 202, 205, 204, 204, 199, 202, 201, 202, 200, 203, 201, 204, 205, 203, 201, 204, 205, 208, 207, 208, 207, 206, 210, 208, 205, 204, 204, 207, 207, 208, 203, 207, 205, 206, 204, 203, 200, 201, 205, 203, 205, 205, 207, 208, 203, 208, 210, 205, 205, 205, 204, 208, 213, 209, 207, 209, 210, 207, 206, 203, 204, 207, 207, 208, 204, 206, 207, 208, 205, 206, 207, 208, 207, 208, 209, 206, 207, 208, 205, 210, 204, 202, 206, 201, 205, 207, 205, 204, 203, 204, 206, 202, 202, 199, 203, 201, 202, 200, 203, 202, 203, 203, 203, 201, 202, 203, 204, 203, 199, 201, 200, 199, 200, 201, 201, 198, 202, 197, 202, 204, 198, 204, 214, 204, 198, 199, 200, 201, 201, 199, 195, 198, 198, 200, 198, 197, 192, 198, 199, 199, 193, 200, 200, 197, 195, 196, 194, 195, 197, 192, 195, 195, 195, 195, 196, 192, 194, 195, 193, 191, 190, 194, 193, 190, 186, 189, 188, 161, 189, 183, 185, 184, 112, 185, 182, 184, 185, 187, 184, 192, 188, 192, 184, 188, 188, 188, 192, 193, 194, 192, 193, 190, 195, 189, 190, 192, 192, 192, 193, 191, 195, 197, 195, 196, 194, 195, 196, 197, 191, 194, 196, 196, 197, 196, 192, 198, 194, 192, 196, 195, 197, 199, 197, 200, 197, 199, 197, 197, 197, 199, 201, 196, 201, 201, 204, 202, 200, 201, 205, 197, 199, 205, 203, 200, 199, 204, 205, 199, 205, 203, 204, 203, 202, 201, 202, 203, 203, 206, 205, 203, 203, 203, 200, 207, 205, 205, 206, 207, 204, 206, 202, 206, 209, 209, 212, 209, 209, 208, 212, 213, 208, 204, 205, 208, 207, 206, 208, 207, 209, 208, 211, 209, 202, 204, 206, 205, 209, 208, 206, 206, 208, 209, 209, 207, 206, 208, 208, 211, 214, 212, 210, 209, 208, 209, 206, 208, 205, 206, 208, 209, 208, 209, 207, 208, 211, 211, 208, 207, 209, 207, 206, 208, 204, 207, 209, 210, 206, 207, 205, 208, 206, 210, 207, 203, 204, 207, 205, 204, 208, 204, 204, 206, 204, 204, 203, 206, 204, 205, 203, 198, 202, 207, 203, 205, 200, 200, 198, 200, 204, 200, 200, 197, 200, 197, 200, 198, 197, 198, 199, 201, 202, 204, 202, 203, 202, 198, 199, 198, 197, 200, 199, 197, 194, 197, 199, 200, 200, 196, 195, 201, 197, 197, 193, 191, 195, 192, 196, 198, 198, 198, 197, 200, 199, 193, 194, 191, 192, 192, 192, 190, 188, 185, 185, 121, 191, 184, 183, 189, 115, 183, 184, 185, 190, 188, 185, 188, 186, 190, 187, 190, 190, 194, 191, 189, 194, 193, 191, 191, 192, 193, 189, 190, 193, 196, 193, 192, 194, 198, 190, 191, 196, 194, 195, 198, 193, 196, 195, 197, 197, 196, 195, 199, 194, 190, 195, 196, 197, 198, 199, 199, 200, 200, 194, 198, 197, 197, 199, 202, 198, 204, 204, 200, 202, 204, 203, 202, 201, 206, 200, 204, 202, 205, 204, 204, 205, 202, 202, 207, 202, 206, 200, 204, 203, 212, 207, 205, 204, 203, 206, 206, 209, 207, 207, 210, 208, 205, 205, 205, 209, 207, 210, 209, 208, 210, 209, 212, 206, 208, 205, 208, 208, 208, 208, 206, 205, 208, 207, 208, 207, 204, 206, 208, 206, 210, 209, 209, 209, 212, 209, 207, 206, 206, 208, 211, 213, 212, 208, 209, 209, 207, 208, 206, 207, 205, 208, 209, 207, 207, 210, 213, 207, 209, 208, 207, 208, 210, 210, 207, 205, 208, 208, 208, 208, 206, 209, 204, 204, 207, 206, 209, 203, 207, 201, 201, 207, 205, 205, 205, 206, 205, 201, 205, 204, 205, 203, 198, 204, 206, 204, 206, 201, 202, 204, 204, 204, 203, 199, 196, 201, 199, 204, 200, 201, 199, 200, 204, 202, 203, 199, 204, 203, 202, 200, 202, 203, 199, 203, 203, 199, 196, 198, 200, 200, 201, 197, 202, 197, 194, 199, 196, 195, 194, 200, 200, 200, 198, 197, 199, 198, 193, 195, 192, 194, 192, 194, 190, 188, 189, 183, 113, 189, 186, 183, 189, 113, 182, 185, 187, 187, 188, 184, 185, 190, 188, 189, 190, 192, 191, 193, 196, 195, 196, 194, 192, 191, 194, 190, 191, 198, 189, 193, 191, 192, 196, 193, 191, 193, 192, 193, 199, 197, 195, 197, 198, 201, 199, 200, 196, 199, 196, 198, 198, 201, 198, 198, 199, 200, 202, 198, 203, 198, 200, 201, 203, 202, 205, 201, 204, 201, 199, 199, 199, 200, 201, 203, 200, 201, 206, 205, 205, 203, 205, 208, 204, 207, 206, 200, 205, 204, 208, 205, 201, 204, 205, 204, 205, 208, 209, 209, 209, 209, 204, 205, 206, 207, 211, 210, 207, 208, 205, 209, 210, 209, 207, 206, 209, 209, 207, 211, 207, 206, 206, 208, 208, 206, 206, 210, 209, 208, 210, 209, 208, 209, 209, 208, 206, 206, 211, 212, 212, 214, 211, 208, 209, 209, 208, 207, 202, 207, 208, 210, 208, 208, 210, 208, 210, 211, 208, 205, 205, 210, 210, 212, 209, 209, 205, 208, 209, 205, 206, 207, 202, 207, 205, 206, 205, 204, 208, 202, 206, 207, 206, 207, 205, 204, 201, 205, 205, 205, 206, 202, 198, 203, 203, 206, 208, 201, 203, 204, 205, 203, 202, 200, 199, 202, 202, 200, 198, 204, 199, 200, 204, 203, 205, 201, 200, 203, 203, 204, 204, 203, 203, 202, 202, 200, 199, 198, 201, 199, 198, 198, 202, 199, 197, 195, 197, 198, 194, 197, 196, 199, 194, 195, 199, 195, 194, 195, 193, 196, 195, 189, 194, 184, 185, 182, 115, 186, 182, 180, 189, 120, 187, 189, 187, 188, 182, 185, 184, 184, 185, 186, 191, 188, 192, 196, 195, 195, 198, 193, 189, 191, 192, 193, 190, 193, 192, 194, 192, 192, 195, 191, 194, 190, 191, 194, 198, 198, 195, 198, 197, 203, 201, 199, 195, 195, 198, 198, 198, 201, 200, 199, 200, 198, 196, 197, 201, 198, 201, 200, 198, 202, 203, 201, 201, 204, 199, 201, 201, 201, 202, 206, 206, 201, 205, 205, 207, 205, 204, 206, 204, 204, 203, 200, 200, 203, 205, 204, 203, 203, 206, 207, 206, 208, 207, 207, 207, 208, 204, 203, 207, 208, 209, 211, 210, 206, 209, 210, 211, 208, 207, 206, 211, 211, 205, 210, 206, 207, 212, 206, 208, 208, 204, 206, 205, 207, 210, 209, 208, 207, 208, 207, 209, 212, 211, 212, 212, 214, 210, 210, 213, 210, 210, 208, 207, 208, 209, 211, 209, 210, 213, 209, 210, 209, 212, 207, 205, 209, 212, 208, 209, 210, 207, 208, 209, 207, 209, 208, 205, 207, 208, 205, 208, 204, 206, 206, 208, 208, 207, 206, 204, 210, 203, 206, 204, 203, 204, 203, 200, 203, 207, 204, 205, 204, 205, 205, 203, 204, 206, 200, 200, 202, 202, 204, 201, 202, 203, 200, 206, 203, 206, 204, 202, 203, 204, 205, 200, 199, 200, 202, 204, 199, 203, 197, 200, 198, 197, 205, 199, 203, 196, 199, 197, 197, 198, 197, 198, 202, 195, 197, 196, 193, 197, 195, 195, 193, 198, 196, 193, 190, 188, 186, 131, 187, 185, 187, 192, 107, 184, 193, 192, 185, 188, 185, 187, 185, 188, 188, 188, 189, 193, 194, 195, 195, 193, 193, 191, 195, 193, 191, 192, 194, 192, 193, 192, 192, 194, 194, 195, 195, 192, 197, 196, 201, 197, 194, 198, 200, 201, 199, 198, 198, 198, 199, 198, 199, 200, 194, 199, 194, 197, 200, 202, 203, 201, 201, 202, 203, 202, 201, 202, 202, 200, 200, 202, 203, 206, 205, 203, 204, 208, 210, 208, 204, 202, 204, 200, 202, 200, 200, 199, 202, 204, 205, 206, 205, 205, 206, 207, 209, 208, 207, 209, 206, 207, 205, 207, 209, 208, 208, 209, 209, 210, 208, 209, 211, 208, 208, 208, 211, 208, 204, 206, 204, 207, 207, 204, 205, 208, 210, 211, 209, 208, 207, 208, 207, 209, 210, 210, 214, 212, 211, 209, 211, 208, 208, 210, 207, 211, 207, 209, 208, 206, 216, 215, 212, 211, 210, 213, 207, 214, 206, 208, 209, 211, 210, 213, 211, 210, 211, 206, 210, 211, 206, 204, 210, 206, 203, 205, 205, 206, 205, 208, 206, 204, 208, 207, 206, 206, 204, 204, 203, 206, 203, 201, 205, 204, 206, 208, 204, 202, 204, 203, 202, 206, 200, 203, 204, 201, 203, 203, 204, 202, 202, 200, 202, 206, 200, 203, 202, 202, 202, 202, 199, 202, 202, 200, 203, 202, 203, 205, 197, 199, 202, 198, 201, 200, 200, 195, 197, 197, 197, 200, 197, 197, 195, 196, 193, 196, 198, 200, 198, 198, 198, 193, 195, 187, 181, 119, 190, 188, 186, 190, 115, 184, 190, 188, 189, 185, 183, 185, 184, 188, 186, 190, 192, 194, 194, 198, 194, 193, 194, 194, 192, 190, 189, 189, 192, 193, 192, 193, 190, 193, 196, 195, 194, 193, 195, 200, 199, 193, 198, 199, 197, 200, 199, 199, 199, 196, 203, 197, 199, 198, 197, 198, 200, 201, 197, 204, 204, 204, 203, 200, 200, 202, 204, 203, 200, 201, 201, 204, 203, 205, 205, 203, 208, 207, 209, 208, 203, 200, 204, 204, 203, 201, 202, 203, 205, 205, 207, 206, 206, 207, 207, 210, 209, 209, 208, 209, 206, 204, 204, 205, 207, 207, 211, 208, 210, 207, 210, 207, 210, 207, 210, 207, 210, 208, 207, 206, 205, 209, 210, 204, 203, 204, 204, 207, 208, 207, 212, 211, 211, 207, 212, 207, 212, 210, 209, 209, 213, 208, 209, 210, 211, 211, 207, 212, 210, 211, 210, 213, 211, 209, 208, 212, 210, 211, 209, 208, 210, 212, 212, 208, 210, 213, 209, 209, 212, 209, 205, 207, 209, 209, 207, 207, 208, 206, 205, 206, 208, 208, 206, 208, 206, 209, 208, 204, 207, 211, 203, 207, 206, 207, 208, 207, 203, 204, 206, 208, 206, 204, 208, 203, 205, 202, 203, 201, 201, 203, 205, 204, 204, 202, 201, 203, 203, 203, 204, 200, 203, 205, 203, 207, 203, 203, 200, 204, 200, 200, 202, 200, 202, 199, 201, 199, 199, 194, 196, 193, 192, 192, 193, 196, 195, 195, 194, 196, 195, 197, 198, 196, 192, 189, 182, 106, 189, 184, 185, 188, 102, 184, 191, 191, 183, 186, 185, 188, 183, 186, 188, 190, 189, 189, 195, 195, 196, 190, 191, 193, 187, 189, 192, 191, 191, 197, 192, 195, 193, 197, 197, 192, 194, 197, 197, 201, 197, 198, 198, 197, 201, 201, 201, 199, 198, 198, 201, 201, 197, 201, 199, 200, 199, 199, 201, 201, 201, 205, 203, 201, 203, 200, 206, 201, 204, 203, 206, 204, 205, 204, 202, 204, 205, 208, 206, 207, 204, 201, 203, 201, 202, 204, 205, 207, 210, 205, 206, 204, 206, 206, 207, 211, 211, 207, 207, 211, 207, 207, 208, 207, 210, 209, 209, 209, 209, 206, 211, 207, 207, 209, 208, 205, 211, 209, 209, 203, 204, 206, 209, 206, 209, 205, 207, 204, 207, 207, 211, 209, 208, 208, 207, 208, 209, 210, 211, 211, 213, 211, 210, 211, 211, 211, 211, 210, 211, 212, 210, 207, 213, 211, 212, 210, 211, 211, 211, 209, 212, 211, 215, 208, 210, 209, 211, 212, 210, 210, 208, 207, 208, 208, 208, 208, 205, 205, 208, 207, 207, 209, 209, 206, 208, 210, 207, 209, 206, 207, 207, 206, 207, 208, 209, 208, 208, 203, 209, 203, 208, 209, 205, 203, 204, 204, 202, 202, 201, 202, 201, 202, 203, 199, 203, 202, 205, 209, 208, 201, 204, 205, 207, 207, 206, 204, 201, 205, 202, 201, 202, 201, 199, 200, 200, 197, 201, 199, 197, 198, 199, 193, 196, 202, 200, 196, 196, 199, 198, 199, 201, 196, 192, 192, 183, 107, 185, 185, 182, 186, 117, 187, 191, 191, 185, 191, 184, 188, 186, 188, 189, 189, 189, 196, 195, 192, 193, 194, 193, 195, 195, 193, 192, 194, 193, 194, 194, 193, 195, 198, 194, 197, 197, 193, 196, 200, 199, 200, 201, 200, 205, 200, 199, 203, 201, 196, 200, 201, 200, 197, 199, 201, 203, 201, 201, 204, 201, 206, 205, 202, 204, 204, 206, 203, 207, 203, 204, 202, 204, 204, 203, 197, 201, 207, 208, 209, 205, 205, 202, 205, 205, 206, 206, 208, 210, 207, 207, 204, 206, 208, 210, 212, 210, 208, 205, 206, 208, 207, 207, 209, 210, 210, 208, 207, 205, 209, 210, 210, 208, 207, 207, 209, 208, 207, 207, 209, 208, 212, 206, 207, 206, 207, 208, 203, 202, 207, 207, 208, 209, 207, 202, 203, 206, 207, 213, 211, 214, 211, 208, 213, 211, 212, 212, 211, 208, 212, 212, 209, 211, 210, 211, 210, 210, 210, 208, 211, 209, 213, 210, 209, 208, 210, 208, 210, 211, 211, 207, 204, 209, 208, 208, 206, 211, 209, 206, 207, 204, 203, 207, 206, 209, 206, 203, 208, 206, 205, 205, 208, 209, 209, 208, 209, 207, 203, 207, 208, 207, 205, 206, 206, 208, 205, 201, 203, 202, 204, 204, 203, 207, 203, 201, 203, 203, 207, 206, 203, 208, 209, 206, 210, 205, 203, 206, 206, 203, 202, 200, 200, 201, 200, 202, 198, 198, 198, 197, 197, 197, 194, 195, 201, 202, 197, 199, 203, 201, 203, 200, 199, 196, 193, 188, 114, 188, 186, 178, 191, 116, 185, 190, 194, 188, 192, 187, 191, 186, 185, 190, 186, 190, 192, 193, 193, 192, 192, 195, 195, 190, 196, 195, 191, 197, 196, 192, 195, 194, 196, 195, 198, 196, 197, 200, 203, 200, 199, 201, 200, 203, 203, 203, 203, 204, 199, 200, 204, 202, 195, 197, 200, 202, 202, 204, 203, 202, 205, 204, 203, 201, 205, 205, 206, 206, 203, 204, 203, 207, 207, 205, 197, 198, 207, 210, 210, 206, 205, 201, 207, 202, 208, 207, 205, 210, 209, 207, 208, 205, 210, 208, 211, 210, 207, 205, 213, 210, 210, 206, 209, 212, 208, 210, 210, 205, 209, 214, 211, 210, 209, 207, 207, 208, 210, 208, 208, 208, 207, 205, 206, 207, 207, 206, 206, 209, 208, 206, 210, 207, 205, 203, 206, 210, 211, 213, 213, 213, 212, 210, 209, 209, 209, 211, 213, 210, 212, 212, 209, 205, 205, 207, 208, 210, 212, 208, 211, 210, 208, 212, 207, 206, 213, 207, 209, 203, 206, 204, 206, 212, 210, 208, 205, 209, 207, 208, 208, 206, 204, 207, 206, 208, 211, 208, 210, 207, 210, 206, 203, 211, 209, 209, 207, 206, 205, 205, 203, 208, 206, 206, 203, 209, 204, 203, 203, 202, 204, 206, 202, 203, 202, 201, 201, 203, 206, 207, 207, 209, 209, 210, 208, 207, 204, 203, 203, 203, 204, 199, 202, 204, 200, 203, 200, 198, 202, 202, 199, 196, 197, 196, 199, 199, 199, 197, 201, 201, 202, 197, 200, 195, 196, 188, 122, 188, 186, 187, 188, 105, 189, 193, 191, 185, 190, 189, 195, 192, 189, 186, 188, 191, 195, 194, 193, 189, 197, 192, 195, 198, 194, 200, 200, 196, 192, 192, 195, 194, 197, 196, 196, 199, 198, 199, 202, 202, 202, 199, 200, 203, 204, 201, 200, 202, 201, 201, 203, 200, 197, 197, 200, 203, 204, 206, 204, 203, 206, 203, 205, 202, 202, 206, 208, 205, 204, 202, 202, 206, 205, 204, 207, 207, 207, 209, 209, 204, 204, 202, 205, 207, 210, 208, 207, 206, 205, 206, 206, 207, 207, 209, 208, 213, 209, 210, 213, 211, 210, 203, 207, 207, 207, 209, 213, 212, 208, 211, 216, 210, 211, 210, 208, 210, 210, 208, 209, 206, 206, 208, 202, 203, 205, 205, 206, 209, 208, 206, 209, 210, 210, 205, 206, 212, 210, 212, 216, 215, 214, 211, 212, 210, 211, 211, 208, 214, 213, 213, 210, 206, 209, 207, 208, 213, 211, 211, 212, 209, 213, 210, 212, 213, 214, 208, 208, 210, 206, 210, 209, 210, 211, 210, 209, 207, 209, 210, 209, 207, 208, 208, 208, 208, 205, 207, 204, 207, 209, 208, 205, 208, 205, 209, 209, 208, 204, 205, 206, 208, 206, 205, 203, 206, 207, 206, 205, 205, 205, 209, 204, 207, 201, 204, 199, 205, 208, 207, 207, 204, 209, 208, 207, 206, 206, 203, 207, 204, 200, 203, 197, 203, 206, 203, 200, 206, 204, 205, 203, 196, 195, 199, 197, 200, 200, 199, 202, 201, 204, 198, 202, 202, 195, 192, 134, 190, 184, 186, 186, 116, 186, 193, 188, 186, 187, 188, 192, 193, 192, 190, 189, 193, 191, 195, 194, 195, 197, 196, 196, 197, 196, 198, 200, 195, 198, 196, 199, 196, 199, 199, 198, 198, 196, 200, 202, 201, 201, 201, 204, 204, 201, 202, 201, 204, 203, 206, 203, 202, 201, 199, 201, 207, 206, 203, 203, 202, 206, 207, 202, 207, 203, 204, 205, 206, 204, 205, 204, 207, 202, 206, 205, 208, 209, 209, 205, 207, 201, 204, 204, 207, 211, 208, 207, 209, 206, 208, 206, 208, 205, 211, 210, 212, 213, 213, 213, 214, 212, 208, 208, 207, 210, 212, 214, 213, 212, 212, 215, 214, 216, 212, 208, 210, 210, 207, 208, 204, 204, 209, 204, 207, 204, 204, 206, 210, 212, 209, 211, 209, 212, 210, 207, 210, 213, 212, 217, 212, 210, 211, 206, 210, 210, 213, 213, 212, 212, 216, 213, 209, 210, 212, 211, 215, 212, 210, 207, 209, 211, 211, 213, 214, 214, 212, 211, 211, 208, 208, 209, 212, 210, 210, 207, 210, 211, 210, 207, 208, 205, 211, 212, 209, 209, 206, 206, 210, 205, 207, 207, 206, 205, 209, 207, 208, 206, 204, 204, 205, 206, 203, 207, 207, 207, 206, 208, 208, 205, 210, 207, 209, 205, 204, 204, 201, 206, 203, 204, 208, 205, 204, 207, 208, 203, 206, 205, 205, 202, 205, 200, 205, 207, 200, 202, 202, 204, 205, 204, 198, 199, 198, 200, 201, 200, 199, 204, 207, 201, 203, 201, 201, 199, 190, 127, 187, 185, 186, 192, 104, 194, 192, 189, 188, 188, 186, 184, 192, 190, 188, 192, 191, 192, 192, 195, 195, 195, 194, 198, 199, 196, 197, 197, 197, 196, 198, 198, 196, 196, 196, 196, 194, 199, 198, 200, 199, 202, 202, 201, 206, 201, 205, 202, 201, 201, 203, 200, 198, 198, 198, 201, 204, 206, 201, 204, 205, 204, 209, 204, 205, 206, 209, 207, 208, 207, 205, 205, 205, 204, 205, 205, 207, 208, 209, 205, 206, 204, 206, 207, 206, 207, 206, 209, 208, 209, 211, 210, 205, 207, 207, 212, 209, 209, 213, 212, 211, 211, 209, 207, 209, 210, 209, 212, 210, 211, 213, 211, 212, 211, 211, 209, 208, 207, 209, 211, 208, 207, 207, 206, 203, 207, 202, 205, 209, 208, 207, 209, 211, 211, 208, 208, 210, 214, 212, 214, 212, 212, 214, 208, 210, 213, 213, 210, 211, 214, 214, 212, 208, 211, 214, 211, 212, 212, 208, 211, 209, 210, 210, 211, 212, 211, 210, 210, 212, 209, 208, 210, 210, 212, 211, 209, 210, 212, 211, 210, 209, 205, 210, 209, 207, 208, 206, 208, 211, 208, 209, 207, 207, 211, 208, 210, 211, 205, 207, 207, 205, 206, 208, 207, 206, 211, 208, 206, 207, 206, 206, 208, 207, 209, 205, 202, 204, 203, 203, 207, 207, 205, 209, 210, 206, 206, 210, 206, 205, 203, 201, 205, 201, 204, 206, 205, 204, 208, 205, 201, 198, 201, 199, 198, 201, 204, 199, 201, 205, 202, 203, 201, 200, 198, 193, 141, 188, 186, 183, 188, 109, 187, 190, 185, 189, 193, 189, 188, 194, 192, 190, 192, 193, 192, 193, 192, 195, 193, 197, 196, 202, 197, 198, 196, 194, 199, 199, 199, 197, 199, 192, 200, 197, 200, 199, 197, 199, 204, 201, 203, 205, 204, 202, 204, 200, 205, 203, 204, 197, 197, 200, 203, 205, 203, 203, 205, 202, 205, 209, 206, 205, 206, 208, 205, 206, 205, 204, 204, 206, 205, 203, 204, 204, 205, 207, 208, 206, 208, 207, 209, 207, 208, 208, 208, 211, 210, 211, 210, 207, 209, 208, 210, 208, 209, 211, 213, 213, 209, 209, 211, 211, 208, 208, 211, 212, 210, 213, 216, 215, 212, 212, 212, 212, 210, 207, 210, 209, 209, 207, 209, 205, 208, 204, 201, 207, 207, 211, 210, 206, 213, 207, 207, 213, 211, 214, 213, 210, 209, 212, 210, 213, 211, 211, 212, 212, 213, 211, 209, 211, 213, 211, 213, 214, 215, 211, 212, 214, 211, 212, 210, 212, 209, 211, 208, 210, 210, 207, 211, 212, 211, 211, 213, 212, 212, 211, 206, 208, 206, 212, 209, 210, 208, 208, 211, 208, 210, 211, 207, 207, 208, 207, 209, 209, 210, 209, 206, 205, 208, 208, 208, 208, 206, 209, 207, 207, 207, 205, 206, 205, 209, 205, 206, 203, 209, 207, 207, 208, 210, 208, 209, 208, 207, 208, 203, 207, 200, 204, 206, 202, 206, 210, 206, 205, 206, 204, 202, 201, 199, 198, 198, 202, 201, 195, 201, 202, 204, 204, 207, 201, 195, 191, 144, 192, 187, 183, 187, 107, 190, 192, 190, 188, 189, 187, 191, 192, 193, 196, 188, 195, 196, 197, 194, 191, 198, 199, 195, 198, 196, 198, 197, 196, 196, 198, 196, 198, 198, 196, 198, 197, 197, 197, 198, 201, 201, 205, 205, 205, 205, 204, 204, 203, 201, 203, 204, 201, 202, 207, 204, 206, 206, 203, 202, 204, 205, 204, 206, 204, 205, 204, 205, 205, 205, 205, 204, 205, 206, 204, 206, 206, 206, 209, 211, 207, 209, 208, 208, 210, 209, 206, 208, 210, 213, 210, 211, 212, 213, 209, 210, 210, 210, 209, 212, 212, 214, 209, 211, 213, 214, 211, 213, 212, 213, 215, 214, 215, 213, 213, 213, 210, 210, 207, 207, 213, 211, 208, 213, 209, 207, 204, 203, 207, 206, 208, 209, 209, 209, 213, 208, 212, 212, 212, 211, 212, 209, 207, 211, 211, 210, 213, 213, 212, 213, 211, 212, 215, 211, 210, 212, 216, 213, 212, 212, 214, 214, 212, 212, 212, 212, 211, 207, 210, 209, 208, 209, 211, 211, 209, 210, 211, 214, 209, 211, 208, 205, 210, 211, 212, 206, 208, 210, 209, 213, 210, 208, 206, 209, 207, 209, 211, 208, 213, 208, 206, 210, 208, 206, 209, 203, 207, 208, 207, 208, 208, 208, 209, 207, 206, 210, 208, 207, 209, 206, 207, 206, 210, 210, 209, 205, 206, 204, 205, 204, 203, 207, 206, 208, 208, 207, 207, 206, 206, 204, 201, 201, 203, 199, 205, 199, 201, 202, 203, 204, 206, 205, 200, 196, 188, 142, 191, 189, 184, 189, 98, 186, 187, 188, 194, 189, 191, 191, 194, 193, 194, 197, 195, 194, 196, 195, 197, 197, 202, 200, 199, 198, 196, 197, 199, 198, 198, 203, 199, 197, 198, 202, 198, 199, 195, 194, 201, 204, 203, 203, 208, 203, 200, 202, 203, 207, 205, 206, 202, 200, 202, 204, 205, 205, 203, 204, 203, 205, 202, 202, 206, 207, 207, 206, 209, 207, 203, 203, 205, 207, 207, 209, 202, 205, 207, 211, 207, 209, 208, 209, 210, 209, 208, 210, 213, 214, 210, 212, 208, 213, 212, 212, 209, 211, 211, 211, 212, 215, 213, 211, 214, 213, 214, 212, 214, 215, 215, 217, 217, 215, 217, 214, 211, 209, 211, 209, 212, 210, 207, 211, 211, 210, 208, 205, 207, 209, 212, 210, 210, 213, 212, 212, 212, 213, 215, 215, 213, 212, 207, 213, 212, 211, 209, 213, 214, 214, 217, 217, 213, 211, 211, 217, 213, 216, 213, 213, 214, 212, 216, 213, 212, 208, 210, 207, 204, 210, 207, 207, 211, 215, 212, 209, 212, 216, 209, 212, 209, 209, 210, 211, 209, 204, 209, 212, 210, 214, 212, 206, 207, 210, 208, 211, 209, 208, 209, 209, 207, 207, 207, 207, 211, 206, 209, 204, 209, 210, 209, 207, 207, 209, 209, 208, 205, 208, 204, 210, 207, 210, 213, 211, 209, 205, 205, 206, 202, 205, 204, 207, 207, 210, 206, 203, 205, 206, 206, 206, 203, 202, 200, 203, 206, 204, 204, 200, 200, 202, 204, 201, 199, 194, 191, 140, 195, 188, 187, 187, 110, 189, 190, 192, 190, 190, 185, 189, 193, 191, 192, 190, 193, 197, 201, 194, 196, 196, 200, 198, 197, 198, 196, 194, 195, 197, 198, 203, 199, 204, 200, 203, 199, 201, 199, 201, 202, 202, 200, 201, 191, 204, 202, 202, 204, 204, 206, 207, 205, 203, 205, 205, 205, 205, 204, 203, 205, 207, 203, 203, 205, 206, 209, 202, 204, 208, 204, 206, 209, 208, 211, 210, 206, 207, 206, 207, 211, 208, 208, 210, 212, 211, 211, 212, 210, 214, 212, 213, 211, 210, 213, 213, 212, 209, 214, 211, 214, 213, 212, 213, 214, 214, 213, 213, 214, 214, 213, 217, 217, 218, 215, 213, 208, 208, 209, 208, 209, 210, 209, 211, 211, 207, 209, 206, 208, 210, 210, 208, 210, 214, 215, 213, 216, 216, 219, 215, 215, 214, 212, 211, 213, 211, 214, 215, 214, 213, 217, 216, 215, 214, 211, 216, 216, 218, 216, 215, 211, 212, 215, 214, 211, 213, 209, 207, 210, 210, 208, 210, 210, 211, 208, 213, 207, 215, 206, 211, 211, 212, 212, 213, 212, 205, 209, 210, 209, 211, 211, 209, 208, 203, 210, 208, 209, 209, 209, 210, 211, 212, 210, 209, 212, 209, 210, 212, 205, 208, 210, 208, 209, 208, 207, 206, 205, 204, 205, 209, 204, 214, 212, 213, 210, 210, 210, 209, 208, 209, 205, 211, 210, 209, 209, 206, 207, 205, 204, 205, 205, 201, 201, 203, 205, 204, 206, 205, 203, 203, 206, 203, 200, 198, 193, 143, 196, 190, 190, 189, 106, 185, 194, 191, 193, 189, 184, 187, 191, 197, 192, 193, 194, 196, 198, 197, 197, 197, 199, 197, 196, 199, 196, 199, 197, 203, 198, 202, 199, 206, 204, 202, 199, 200, 198, 198, 201, 202, 202, 201, 200, 205, 204, 205, 208, 203, 208, 204, 205, 202, 208, 206, 206, 206, 203, 205, 206, 209, 208, 205, 205, 203, 209, 205, 208, 208, 208, 209, 212, 210, 213, 210, 208, 208, 208, 207, 211, 206, 208, 210, 212, 214, 209, 212, 212, 211, 210, 211, 210, 211, 213, 210, 211, 213, 215, 215, 213, 212, 213, 214, 213, 214, 214, 212, 214, 213, 214, 216, 217, 216, 214, 214, 211, 208, 209, 209, 209, 210, 212, 211, 212, 210, 211, 209, 209, 210, 211, 209, 210, 212, 214, 215, 214, 212, 216, 213, 216, 213, 210, 214, 211, 213, 213, 214, 214, 215, 216, 218, 216, 212, 212, 209, 217, 214, 214, 212, 214, 215, 212, 212, 213, 211, 211, 208, 209, 213, 210, 211, 214, 208, 209, 212, 212, 213, 213, 210, 209, 210, 210, 211, 209, 208, 204, 204, 209, 211, 207, 207, 210, 208, 212, 213, 208, 212, 209, 207, 209, 209, 210, 210, 210, 212, 211, 209, 207, 207, 208, 208, 208, 207, 207, 207, 204, 207, 204, 205, 207, 212, 210, 214, 210, 210, 212, 212, 209, 208, 209, 208, 210, 209, 211, 209, 207, 204, 206, 205, 208, 203, 203, 204, 206, 209, 205, 206, 204, 204, 207, 203, 200, 196, 191, 139, 195, 189, 191, 190, 106, 189, 192, 190, 190, 189, 193, 196, 194, 195, 190, 194, 196, 201, 198, 195, 196, 196, 196, 198, 198, 195, 198, 197, 195, 199, 200, 202, 200, 204, 203, 201, 200, 202, 199, 202, 203, 202, 202, 205, 207, 207, 208, 211, 207, 207, 207, 205, 207, 204, 206, 208, 206, 205, 205, 206, 208, 207, 206, 209, 208, 211, 213, 211, 212, 208, 210, 210, 212, 211, 213, 208, 210, 209, 210, 211, 209, 211, 211, 212, 211, 211, 211, 212, 212, 213, 205, 212, 211, 212, 211, 212, 213, 213, 213, 215, 213, 210, 212, 215, 214, 213, 214, 214, 213, 212, 214, 216, 215, 216, 211, 213, 212, 209, 212, 209, 212, 210, 216, 214, 213, 213, 210, 210, 211, 211, 206, 212, 212, 213, 217, 216, 214, 216, 219, 217, 213, 214, 214, 216, 212, 214, 216, 213, 215, 219, 218, 217, 216, 209, 212, 212, 215, 214, 216, 215, 214, 217, 214, 214, 211, 212, 211, 211, 214, 212, 212, 211, 213, 210, 213, 211, 210, 211, 215, 214, 211, 209, 211, 209, 210, 205, 206, 206, 210, 210, 214, 209, 209, 207, 210, 211, 208, 208, 210, 210, 210, 212, 211, 213, 211, 213, 210, 207, 209, 211, 209, 209, 206, 211, 206, 207, 208, 205, 211, 209, 205, 211, 214, 212, 211, 211, 211, 212, 211, 212, 211, 211, 209, 214, 212, 212, 208, 204, 206, 207, 207, 205, 205, 208, 207, 207, 210, 208, 206, 210, 206, 201, 197, 202, 192, 138, 192, 190, 187, 191, 116, 189, 195, 193, 192, 191, 194, 194, 192, 198, 198, 196, 197, 199, 202, 201, 198, 197, 197, 200, 200, 197, 199, 197, 199, 199, 200, 202, 206, 202, 202, 204, 202, 202, 200, 198, 203, 202, 205, 203, 205, 205, 209, 207, 206, 205, 207, 206, 208, 207, 207, 208, 206, 204, 206, 204, 208, 206, 207, 209, 207, 210, 211, 214, 215, 212, 210, 208, 213, 213, 211, 209, 211, 208, 209, 213, 211, 212, 212, 212, 214, 209, 211, 212, 214, 216, 213, 211, 214, 211, 214, 216, 215, 213, 215, 213, 213, 213, 215, 215, 217, 213, 215, 213, 212, 214, 214, 218, 216, 216, 214, 214, 215, 211, 213, 209, 210, 214, 216, 214, 216, 214, 212, 211, 212, 212, 212, 215, 211, 213, 216, 215, 218, 216, 216, 216, 215, 214, 213, 216, 213, 213, 216, 216, 216, 217, 215, 214, 215, 214, 213, 216, 217, 215, 214, 210, 212, 212, 214, 213, 210, 212, 212, 213, 218, 214, 210, 216, 213, 213, 212, 209, 215, 213, 213, 215, 210, 209, 214, 209, 210, 204, 205, 206, 212, 210, 210, 211, 209, 205, 212, 212, 210, 207, 210, 211, 215, 212, 213, 212, 214, 214, 209, 207, 211, 210, 209, 212, 208, 209, 213, 207, 210, 211, 210, 209, 212, 214, 215, 215, 211, 210, 212, 212, 213, 214, 213, 211, 211, 209, 210, 209, 207, 210, 209, 213, 207, 207, 208, 207, 209, 207, 208, 211, 208, 209, 211, 205, 202, 198, 191, 145, 195, 195, 189, 196, 116, 192, 193, 196, 193, 197, 198, 197, 198, 197, 199, 194, 197, 199, 205, 199, 200, 201, 202, 201, 201, 198, 201, 201, 199, 199, 200, 202, 201, 203, 202, 208, 203, 205, 203, 202, 204, 201, 206, 203, 208, 206, 206, 208, 209, 208, 210, 210, 209, 203, 209, 207, 207, 207, 206, 207, 209, 204, 210, 208, 212, 211, 212, 213, 213, 213, 210, 209, 210, 210, 212, 211, 207, 210, 211, 214, 213, 209, 209, 212, 217, 211, 212, 213, 215, 216, 212, 208, 212, 210, 212, 214, 216, 212, 211, 214, 213, 212, 213, 212, 212, 211, 214, 214, 210, 214, 218, 217, 216, 217, 217, 214, 212, 210, 212, 209, 212, 213, 215, 213, 215, 213, 213, 211, 210, 211, 213, 212, 212, 214, 217, 214, 217, 216, 216, 215, 213, 213, 215, 215, 218, 214, 216, 214, 214, 215, 219, 218, 215, 216, 217, 215, 219, 214, 214, 213, 215, 212, 213, 214, 214, 216, 215, 215, 220, 217, 215, 214, 217, 214, 211, 211, 213, 212, 215, 213, 210, 208, 212, 210, 211, 205, 204, 208, 212, 212, 208, 212, 212, 209, 212, 211, 208, 208, 210, 210, 213, 213, 215, 214, 216, 213, 210, 210, 209, 211, 208, 211, 209, 207, 211, 209, 210, 207, 208, 210, 214, 214, 218, 215, 213, 215, 215, 215, 215, 215, 213, 210, 211, 213, 215, 210, 205, 210, 209, 213, 208, 208, 211, 211, 213, 215, 209, 208, 209, 207, 210, 207, 203, 200, 198, 150, 194, 195, 189, 195, 130, 192, 199, 192, 192, 197, 195, 195, 197, 194, 198, 196, 197, 201, 197, 201, 201, 196, 201, 203, 202, 201, 198, 197, 196, 198, 203, 205, 206, 207, 204, 204, 205, 205, 204, 205, 206, 204, 206, 203, 207, 209, 208, 206, 208, 208, 209, 209, 209, 205, 208, 211, 205, 210, 209, 209, 210, 208, 211, 210, 211, 209, 212, 212, 214, 213, 208, 212, 209, 212, 212, 216, 210, 215, 214, 213, 212, 210, 212, 213, 211, 210, 210, 212, 213, 211, 204, 210, 212, 213, 214, 213, 213, 213, 211, 216, 213, 214, 214, 213, 213, 212, 214, 211, 212, 216, 215, 219, 217, 218, 218, 214, 214, 211, 212, 213, 213, 212, 215, 213, 214, 211, 212, 214, 212, 213, 212, 211, 214, 216, 218, 216, 217, 216, 214, 215, 215, 217, 217, 217, 215, 216, 216, 217, 216, 217, 219, 217, 215, 214, 215, 215, 217, 216, 215, 218, 215, 214, 213, 217, 218, 216, 216, 217, 215, 217, 214, 216, 217, 217, 214, 212, 213, 214, 216, 215, 212, 213, 211, 213, 212, 207, 206, 212, 213, 212, 212, 213, 211, 211, 213, 214, 211, 209, 209, 213, 216, 216, 213, 213, 216, 213, 212, 211, 208, 214, 208, 211, 211, 209, 214, 208, 214, 215, 210, 213, 217, 214, 214, 215, 213, 214, 216, 214, 216, 214, 213, 217, 214, 214, 210, 211, 209, 210, 210, 214, 211, 210, 211, 209, 212, 217, 209, 212, 209, 207, 207, 207, 206, 202, 198, 161, 195, 195, 189, 192, 115, 195, 194, 194, 196, 201, 196, 200, 195, 195, 199, 200, 198, 202, 201, 199, 200, 200, 202, 200, 201, 204, 201, 200, 200, 200, 203, 207, 206, 206, 205, 201, 207, 207, 206, 206, 207, 202, 202, 203, 204, 206, 208, 209, 209, 209, 210, 213, 209, 205, 208, 207, 204, 208, 209, 208, 212, 211, 212, 213, 210, 211, 212, 213, 214, 214, 210, 211, 212, 214, 214, 216, 212, 214, 212, 211, 211, 210, 212, 212, 213, 213, 210, 209, 213, 216, 209, 213, 216, 215, 213, 216, 214, 209, 209, 214, 216, 212, 213, 212, 214, 215, 214, 212, 215, 215, 214, 218, 217, 216, 217, 217, 214, 209, 213, 214, 212, 210, 213, 212, 212, 211, 213, 215, 211, 213, 216, 214, 215, 216, 219, 217, 216, 212, 217, 214, 216, 216, 216, 217, 217, 218, 215, 214, 217, 218, 217, 218, 217, 218, 215, 218, 217, 216, 215, 215, 214, 216, 218, 219, 219, 218, 215, 217, 215, 214, 213, 215, 218, 215, 216, 215, 214, 216, 218, 218, 211, 213, 216, 218, 216, 213, 213, 209, 215, 213, 215, 212, 215, 213, 216, 214, 212, 211, 213, 212, 213, 215, 213, 216, 215, 211, 214, 210, 209, 211, 213, 213, 212, 213, 216, 214, 212, 213, 215, 214, 216, 216, 219, 214, 212, 215, 213, 215, 215, 211, 214, 215, 215, 214, 211, 213, 208, 208, 212, 207, 214, 209, 208, 211, 208, 207, 209, 210, 206, 208, 207, 206, 211, 204, 198, 175, 198, 190, 189, 191, 124, 192, 197, 195, 194, 199, 200, 197, 194, 195, 197, 201, 197, 199, 200, 198, 202, 198, 205, 203, 205, 203, 203, 204, 203, 201, 202, 203, 202, 203, 205, 205, 204, 207, 204, 206, 205, 204, 204, 204, 206, 205, 211, 207, 207, 210, 212, 213, 209, 210, 209, 211, 208, 208, 208, 206, 209, 209, 210, 209, 209, 210, 212, 211, 210, 212, 210, 210, 209, 214, 213, 212, 213, 211, 214, 213, 213, 209, 209, 213, 214, 213, 215, 212, 215, 216, 215, 216, 214, 214, 215, 213, 215, 213, 214, 215, 214, 217, 216, 217, 217, 214, 216, 212, 212, 214, 213, 215, 214, 216, 214, 214, 218, 211, 214, 214, 214, 212, 213, 212, 210, 213, 215, 211, 214, 215, 214, 216, 215, 216, 219, 216, 216, 215, 215, 216, 217, 220, 216, 215, 220, 220, 216, 216, 218, 217, 218, 219, 217, 217, 217, 218, 220, 217, 219, 216, 215, 218, 218, 219, 219, 218, 220, 218, 214, 213, 213, 215, 218, 220, 217, 214, 212, 210, 216, 216, 210, 214, 214, 216, 214, 214, 214, 212, 212, 213, 215, 212, 213, 216, 214, 212, 209, 209, 213, 215, 212, 216, 209, 216, 216, 213, 213, 213, 211, 212, 210, 212, 213, 210, 214, 214, 213, 216, 217, 214, 215, 214, 217, 213, 212, 211, 212, 215, 213, 213, 213, 213, 212, 211, 210, 212, 211, 208, 212, 213, 213, 212, 212, 210, 207, 209, 210, 207, 207, 210, 209, 209, 206, 205, 196, 166, 195, 190, 191, 196, 132, 195, 197, 198, 197, 197, 198, 198, 197, 196, 197, 198, 203, 202, 201, 199, 199, 200, 200, 203, 200, 199, 200, 200, 200, 200, 206, 203, 202, 202, 206, 209, 207, 205, 206, 205, 205, 205, 207, 209, 209, 209, 210, 208, 209, 213, 214, 209, 212, 208, 210, 211, 212, 211, 212, 209, 208, 212, 213, 213, 212, 211, 209, 208, 210, 209, 208, 211, 212, 214, 212, 215, 215, 212, 214, 213, 212, 210, 210, 214, 212, 213, 212, 215, 214, 216, 214, 214, 214, 217, 219, 216, 215, 213, 213, 213, 216, 216, 213, 217, 216, 217, 218, 214, 214, 216, 214, 216, 218, 218, 216, 214, 213, 215, 212, 213, 211, 210, 212, 210, 210, 214, 213, 214, 216, 214, 213, 216, 218, 218, 216, 216, 216, 215, 217, 217, 218, 218, 220, 219, 221, 222, 220, 218, 217, 218, 219, 218, 217, 216, 217, 216, 220, 218, 215, 215, 218, 217, 218, 218, 219, 217, 217, 216, 216, 214, 215, 212, 217, 215, 215, 212, 211, 212, 215, 214, 215, 216, 219, 214, 217, 214, 212, 215, 216, 212, 210, 216, 214, 216, 214, 212, 212, 213, 211, 219, 212, 213, 212, 217, 216, 216, 213, 216, 213, 211, 213, 217, 216, 211, 213, 214, 213, 214, 217, 218, 216, 214, 215, 217, 212, 211, 214, 212, 215, 214, 216, 214, 214, 210, 209, 212, 212, 214, 214, 214, 213, 213, 214, 210, 211, 208, 210, 207, 210, 209, 212, 211, 206, 207, 199, 156, 193, 191, 193, 198, 134, 190, 196, 198, 193, 198, 198, 199, 199, 200, 200, 200, 200, 201, 203, 202, 199, 201, 202, 204, 199, 202, 202, 202, 199, 204, 206, 205, 203, 206, 204, 207, 204, 206, 205, 205, 205, 205, 207, 207, 214, 210, 212, 208, 210, 213, 211, 210, 214, 210, 212, 212, 212, 211, 207, 208, 210, 208, 215, 213, 211, 213, 213, 213, 211, 211, 211, 209, 214, 215, 214, 214, 216, 214, 214, 213, 212, 211, 212, 215, 214, 212, 208, 215, 215, 216, 219, 214, 216, 216, 218, 219, 216, 215, 214, 218, 217, 218, 218, 220, 218, 218, 216, 217, 216, 213, 216, 218, 218, 216, 217, 214, 217, 217, 215, 214, 212, 210, 215, 214, 216, 215, 215, 215, 216, 214, 210, 216, 217, 216, 216, 216, 216, 214, 215, 216, 221, 219, 219, 218, 223, 221, 223, 219, 217, 219, 218, 219, 216, 217, 216, 221, 220, 217, 213, 216, 220, 218, 217, 216, 217, 218, 220, 220, 218, 215, 216, 216, 218, 218, 218, 213, 212, 213, 216, 216, 216, 210, 214, 217, 218, 213, 210, 214, 213, 213, 215, 215, 215, 216, 215, 216, 216, 217, 213, 216, 211, 213, 213, 212, 215, 214, 215, 215, 217, 216, 212, 212, 217, 214, 214, 214, 212, 215, 219, 216, 215, 218, 219, 216, 215, 214, 213, 213, 214, 218, 215, 215, 212, 212, 215, 215, 217, 214, 217, 214, 212, 214, 212, 211, 213, 208, 209, 208, 209, 209, 211, 210, 208, 205, 197, 145, 195, 195, 192, 197, 121, 194, 194, 193, 198, 196, 198, 201, 200, 196, 197, 193, 195, 203, 199, 203, 199, 201, 203, 204, 203, 204, 201, 201, 201, 203, 206, 201, 203, 205, 205, 209, 204, 208, 205, 206, 205, 207, 206, 210, 210, 211, 213, 211, 210, 213, 213, 213, 213, 208, 212, 212, 211, 212, 211, 206, 212, 213, 218, 208, 211, 212, 216, 215, 210, 213, 214, 214, 212, 215, 214, 213, 212, 214, 212, 212, 209, 213, 208, 214, 211, 213, 214, 214, 215, 219, 217, 214, 218, 217, 218, 217, 217, 216, 213, 215, 216, 215, 217, 217, 215, 216, 217, 217, 219, 216, 219, 218, 218, 216, 213, 218, 215, 215, 215, 213, 212, 216, 215, 216, 213, 216, 216, 218, 215, 215, 215, 217, 218, 217, 217, 215, 216, 213, 216, 218, 220, 219, 218, 218, 221, 221, 221, 219, 221, 220, 218, 220, 216, 218, 218, 218, 218, 218, 217, 216, 219, 218, 219, 219, 219, 216, 218, 217, 215, 216, 221, 216, 219, 218, 218, 214, 210, 216, 214, 217, 213, 212, 215, 217, 214, 213, 213, 215, 216, 214, 215, 214, 212, 219, 215, 213, 215, 218, 218, 216, 210, 217, 215, 214, 213, 213, 214, 215, 215, 216, 218, 214, 214, 214, 212, 214, 219, 216, 219, 218, 216, 217, 217, 216, 215, 214, 213, 213, 217, 216, 211, 214, 216, 217, 216, 215, 216, 212, 217, 213, 215, 215, 211, 213, 213, 212, 209, 211, 209, 210, 212, 211, 208, 205, 197, 145, 196, 194, 192, 198, 117, 195, 199, 197, 198, 198, 198, 201, 197, 196, 195, 197, 198, 202, 201, 202, 200, 198, 206, 203, 205, 206, 203, 204, 204, 203, 206, 204, 204, 204, 206, 206, 207, 207, 205, 207, 206, 206, 211, 210, 212, 211, 213, 211, 210, 211, 210, 211, 212, 208, 209, 216, 210, 207, 211, 210, 210, 213, 216, 213, 213, 213, 216, 218, 215, 213, 212, 214, 215, 214, 215, 212, 210, 213, 216, 212, 212, 212, 210, 212, 213, 213, 215, 215, 217, 217, 217, 215, 217, 213, 215, 220, 218, 216, 215, 214, 216, 219, 214, 217, 219, 218, 217, 217, 217, 217, 216, 216, 217, 216, 218, 218, 217, 217, 215, 216, 215, 216, 215, 216, 214, 219, 217, 216, 217, 220, 217, 218, 217, 216, 215, 215, 217, 213, 218, 221, 220, 218, 220, 220, 220, 221, 220, 218, 219, 218, 218, 217, 217, 217, 221, 221, 218, 218, 216, 218, 219, 219, 220, 216, 216, 217, 216, 217, 216, 218, 219, 219, 219, 220, 217, 216, 216, 217, 218, 214, 210, 212, 213, 216, 214, 214, 217, 214, 217, 216, 216, 216, 217, 215, 219, 215, 215, 214, 215, 217, 215, 213, 216, 214, 214, 215, 212, 216, 215, 215, 218, 217, 217, 213, 213, 212, 213, 214, 218, 217, 215, 219, 218, 217, 215, 217, 216, 216, 214, 216, 213, 214, 217, 216, 216, 215, 215, 215, 214, 217, 218, 215, 213, 213, 213, 214, 209, 210, 210, 213, 214, 211, 209, 205, 199, 150, 199, 197, 194, 199, 126, 195, 201, 200, 195, 200, 196, 201, 203, 196, 201, 198, 195, 201, 198, 199, 204, 203, 208, 204, 205, 206, 204, 205, 205, 202, 205, 205, 208, 204, 209, 207, 207, 207, 206, 206, 208, 206, 206, 208, 210, 210, 211, 211, 209, 208, 211, 210, 211, 209, 212, 213, 209, 213, 211, 213, 212, 213, 215, 212, 212, 211, 215, 214, 211, 211, 212, 215, 217, 213, 215, 214, 209, 214, 214, 215, 213, 212, 211, 215, 211, 216, 214, 216, 216, 218, 216, 217, 215, 214, 218, 220, 216, 213, 217, 218, 213, 218, 218, 216, 220, 219, 220, 219, 217, 214, 217, 218, 217, 216, 217, 216, 218, 219, 217, 217, 216, 217, 215, 218, 218, 217, 214, 213, 215, 217, 217, 215, 215, 216, 219, 216, 221, 216, 217, 220, 223, 219, 220, 220, 221, 222, 221, 220, 220, 218, 219, 221, 219, 216, 220, 218, 219, 220, 217, 220, 219, 219, 218, 215, 216, 216, 216, 216, 214, 219, 219, 218, 221, 220, 217, 216, 214, 217, 216, 211, 213, 214, 217, 218, 213, 215, 213, 214, 218, 217, 217, 216, 218, 217, 217, 216, 218, 213, 216, 217, 216, 217, 215, 217, 217, 216, 216, 217, 217, 217, 217, 219, 216, 214, 212, 211, 213, 215, 215, 216, 214, 218, 217, 216, 217, 214, 216, 217, 217, 215, 218, 215, 217, 216, 218, 215, 213, 215, 214, 217, 217, 217, 213, 214, 212, 214, 211, 212, 211, 212, 216, 214, 207, 205, 201, 159, 198, 193, 192, 201, 124, 192, 199, 197, 196, 196, 200, 200, 200, 196, 198, 195, 197, 207, 204, 207, 201, 206, 207, 205, 210, 207, 210, 207, 210, 206, 204, 208, 206, 205, 207, 207, 208, 206, 208, 205, 206, 206, 207, 211, 210, 212, 213, 211, 210, 212, 214, 214, 213, 211, 214, 213, 210, 213, 211, 214, 215, 214, 214, 214, 215, 212, 214, 213, 213, 214, 217, 214, 216, 214, 212, 212, 213, 214, 218, 219, 212, 212, 211, 215, 214, 213, 216, 212, 216, 220, 220, 219, 216, 216, 218, 221, 216, 213, 215, 216, 216, 220, 221, 219, 218, 220, 218, 217, 218, 214, 217, 218, 216, 221, 216, 215, 217, 216, 215, 217, 216, 217, 216, 216, 215, 216, 218, 215, 215, 218, 216, 217, 216, 215, 217, 217, 217, 217, 218, 222, 221, 218, 222, 221, 221, 221, 222, 222, 220, 220, 220, 219, 221, 217, 218, 221, 220, 217, 217, 218, 217, 220, 218, 217, 218, 215, 221, 221, 219, 220, 217, 221, 221, 218, 214, 216, 220, 216, 218, 215, 215, 213, 218, 217, 215, 215, 214, 212, 216, 216, 217, 219, 219, 219, 221, 218, 216, 215, 215, 218, 218, 218, 216, 215, 216, 217, 218, 215, 216, 217, 219, 219, 214, 214, 215, 216, 218, 217, 218, 217, 219, 221, 219, 215, 216, 215, 218, 217, 217, 216, 215, 213, 214, 217, 216, 214, 213, 213, 215, 214, 212, 216, 213, 210, 212, 216, 208, 210, 211, 215, 216, 213, 211, 208, 198, 155, 202, 193, 195, 196, 117, 193, 201, 198, 196, 196, 202, 198, 201, 199, 197, 198, 197, 199, 206, 205, 209, 206, 209, 208, 209, 209, 209, 206, 210, 202, 203, 208, 203, 204, 206, 206, 205, 205, 206, 208, 209, 206, 211, 212, 215, 214, 213, 211, 210, 213, 216, 213, 211, 211, 214, 215, 213, 213, 216, 217, 217, 215, 218, 214, 216, 212, 213, 216, 214, 216, 216, 216, 214, 216, 210, 212, 212, 213, 217, 217, 215, 213, 215, 216, 213, 211, 214, 215, 216, 217, 218, 217, 214, 215, 221, 217, 217, 217, 214, 218, 217, 218, 220, 216, 219, 220, 219, 217, 216, 217, 219, 218, 218, 220, 219, 216, 220, 219, 218, 220, 219, 216, 217, 216, 215, 216, 219, 218, 218, 219, 216, 217, 212, 218, 219, 215, 216, 217, 223, 223, 223, 221, 222, 222, 224, 221, 221, 223, 222, 222, 218, 219, 217, 216, 218, 222, 218, 218, 217, 221, 219, 220, 218, 217, 214, 221, 221, 221, 222, 219, 221, 223, 222, 218, 218, 217, 218, 219, 218, 215, 214, 215, 215, 218, 218, 215, 216, 216, 218, 219, 218, 218, 218, 219, 219, 219, 217, 219, 215, 216, 219, 217, 222, 215, 217, 219, 219, 218, 216, 216, 221, 219, 218, 214, 216, 216, 218, 217, 217, 216, 221, 220, 220, 216, 216, 213, 216, 220, 216, 217, 219, 218, 215, 218, 219, 217, 217, 214, 217, 217, 215, 215, 214, 213, 213, 213, 213, 209, 212, 215, 213, 215, 211, 204, 198, 159, 202, 196, 192, 199, 103, 189, 198, 197, 197, 198, 195, 201, 199, 198, 195, 198, 197, 199, 205, 202, 205, 207, 208, 207, 208, 206, 205, 204, 207, 202, 202, 203, 205, 207, 205, 208, 208, 205, 204, 210, 212, 209, 213, 210, 212, 213, 210, 211, 207, 214, 214, 213, 214, 213, 217, 216, 217, 215, 214, 215, 218, 217, 219, 216, 212, 213, 214, 217, 216, 214, 218, 219, 216, 214, 214, 210, 212, 214, 215, 214, 215, 215, 215, 215, 215, 214, 217, 214, 217, 216, 219, 221, 217, 217, 220, 220, 216, 214, 217, 220, 220, 218, 219, 216, 220, 219, 218, 218, 216, 218, 220, 217, 219, 217, 217, 218, 218, 218, 219, 218, 218, 215, 215, 216, 217, 216, 217, 219, 215, 218, 215, 214, 216, 219, 219, 218, 219, 219, 222, 222, 222, 223, 222, 221, 223, 220, 219, 220, 221, 220, 218, 218, 218, 218, 219, 223, 223, 218, 218, 221, 220, 221, 218, 216, 218, 219, 220, 219, 218, 218, 219, 224, 223, 220, 217, 216, 217, 217, 217, 217, 214, 215, 216, 216, 215, 217, 216, 219, 217, 218, 216, 216, 220, 218, 219, 216, 212, 216, 216, 219, 217, 218, 215, 214, 218, 216, 216, 219, 216, 215, 218, 216, 215, 220, 216, 216, 218, 216, 217, 217, 217, 219, 219, 218, 218, 215, 216, 219, 221, 217, 216, 214, 218, 216, 216, 215, 215, 216, 212, 214, 214, 212, 215, 215, 214, 216, 211, 213, 209, 213, 216, 216, 212, 207, 196, 151, 199, 196, 195, 198, 115, 193, 199, 194, 194, 196, 198, 202, 199, 197, 198, 201, 201, 203, 203, 205, 206, 205, 206, 205, 208, 203, 207, 208, 206, 205, 210, 205, 205, 204, 207, 210, 209, 209, 205, 211, 209, 210, 210, 214, 212, 212, 209, 208, 208, 214, 215, 212, 214, 214, 214, 212, 216, 214, 218, 216, 216, 216, 219, 212, 212, 215, 216, 217, 214, 217, 219, 221, 219, 216, 218, 212, 209, 213, 214, 215, 216, 214, 214, 215, 216, 217, 216, 215, 218, 218, 218, 220, 221, 216, 221, 218, 218, 217, 214, 219, 219, 220, 219, 218, 218, 220, 218, 220, 217, 215, 217, 219, 218, 218, 218, 218, 218, 218, 221, 219, 218, 215, 218, 215, 215, 218, 218, 217, 220, 217, 218, 217, 218, 218, 216, 220, 219, 218, 220, 221, 225, 221, 222, 221, 222, 221, 220, 220, 222, 220, 222, 221, 217, 219, 222, 220, 221, 223, 223, 218, 220, 223, 221, 216, 218, 218, 220, 222, 219, 220, 221, 224, 223, 223, 221, 217, 218, 218, 218, 217, 211, 216, 216, 216, 215, 213, 218, 219, 220, 220, 216, 216, 218, 219, 219, 218, 217, 217, 216, 218, 217, 222, 218, 217, 220, 218, 218, 218, 217, 216, 218, 216, 214, 219, 215, 215, 218, 219, 216, 217, 217, 219, 219, 217, 218, 217, 217, 220, 221, 220, 217, 217, 220, 215, 217, 217, 213, 213, 213, 218, 217, 215, 212, 214, 215, 217, 211, 214, 208, 215, 213, 213, 213, 209, 203, 156, 198, 198, 195, 198, 103, 192, 194, 196, 192, 201, 199, 202, 198, 198, 203, 197, 202, 202, 202, 206, 208, 207, 209, 207, 204, 205, 206, 206, 211, 209, 213, 208, 206, 207, 209, 209, 207, 208, 209, 211, 213, 211, 211, 209, 211, 212, 209, 210, 209, 213, 216, 211, 214, 213, 218, 214, 217, 215, 217, 214, 217, 216, 217, 212, 216, 215, 218, 216, 215, 217, 217, 219, 217, 220, 215, 217, 213, 217, 215, 216, 216, 217, 216, 217, 217, 216, 216, 215, 219, 219, 219, 220, 219, 216, 219, 220, 218, 217, 217, 219, 220, 219, 220, 219, 219, 222, 219, 219, 215, 216, 218, 216, 220, 219, 221, 218, 219, 219, 219, 216, 217, 216, 218, 218, 218, 215, 219, 216, 218, 216, 218, 219, 219, 220, 219, 220, 221, 221, 218, 221, 223, 219, 221, 223, 223, 220, 221, 222, 222, 223, 222, 218, 218, 218, 222, 222, 223, 223, 222, 220, 220, 222, 221, 218, 218, 218, 220, 223, 222, 219, 222, 223, 221, 224, 220, 218, 221, 219, 219, 219, 214, 216, 216, 217, 216, 213, 221, 216, 217, 215, 217, 218, 218, 218, 218, 219, 218, 216, 220, 218, 221, 219, 220, 219, 220, 218, 218, 221, 216, 216, 216, 215, 219, 219, 218, 215, 216, 217, 219, 215, 218, 217, 218, 219, 217, 216, 216, 221, 217, 222, 218, 218, 220, 216, 218, 213, 214, 210, 219, 216, 213, 217, 215, 217, 216, 215, 214, 213, 213, 215, 217, 216, 210, 210, 202, 154, 202, 194, 197, 197, 91, 192, 197, 196, 198, 200, 198, 200, 202, 201, 198, 201, 202, 204, 205, 206, 208, 209, 208, 208, 206, 205, 208, 207, 211, 209, 211, 208, 211, 209, 210, 208, 206, 209, 212, 210, 212, 212, 214, 210, 212, 213, 211, 209, 212, 212, 216, 216, 217, 216, 216, 215, 217, 217, 213, 217, 219, 216, 218, 216, 216, 217, 216, 219, 214, 216, 216, 217, 217, 216, 216, 218, 215, 216, 218, 217, 217, 219, 216, 220, 216, 217, 218, 217, 219, 216, 219, 220, 218, 216, 218, 219, 221, 218, 218, 219, 220, 217, 222, 222, 220, 222, 220, 218, 215, 216, 221, 220, 223, 223, 220, 217, 220, 221, 221, 218, 216, 215, 221, 219, 219, 214, 220, 216, 216, 218, 218, 218, 217, 218, 220, 219, 222, 220, 222, 220, 223, 220, 222, 224, 223, 222, 224, 221, 221, 223, 221, 221, 219, 221, 220, 223, 222, 223, 219, 222, 224, 225, 222, 219, 222, 220, 218, 223, 221, 219, 218, 221, 221, 220, 219, 219, 221, 220, 219, 220, 216, 217, 220, 218, 218, 217, 221, 218, 220, 213, 219, 218, 219, 218, 217, 219, 213, 217, 220, 218, 220, 220, 221, 221, 219, 216, 221, 221, 217, 214, 216, 215, 218, 219, 220, 215, 218, 219, 221, 216, 216, 217, 217, 220, 217, 216, 219, 220, 223, 221, 219, 218, 217, 215, 214, 213, 211, 213, 215, 218, 217, 219, 217, 218, 217, 217, 212, 213, 214, 212, 216, 214, 213, 208, 201, 156, 200, 198, 195, 198, 89, 190, 198, 196, 196, 198, 201, 200, 201, 203, 200, 203, 207, 208, 206, 207, 205, 206, 211, 203, 210, 210, 210, 210, 211, 210, 209, 209, 210, 211, 210, 210, 207, 210, 212, 211, 212, 214, 212, 212, 211, 211, 213, 213, 212, 213, 213, 217, 217, 217, 216, 216, 218, 216, 214, 218, 217, 217, 219, 217, 216, 217, 218, 219, 215, 218, 215, 216, 216, 220, 216, 217, 216, 216, 220, 217, 219, 218, 218, 219, 216, 218, 216, 217, 218, 217, 219, 217, 218, 216, 218, 220, 217, 220, 218, 219, 220, 221, 221, 222, 219, 219, 219, 220, 216, 220, 220, 221, 218, 221, 221, 221, 221, 223, 220, 218, 217, 217, 221, 220, 219, 217, 218, 217, 218, 219, 217, 219, 218, 218, 218, 218, 221, 222, 220, 222, 222, 224, 222, 224, 223, 222, 224, 220, 219, 223, 219, 220, 221, 219, 220, 224, 223, 221, 219, 223, 224, 222, 222, 220, 219, 220, 218, 222, 221, 219, 219, 220, 221, 222, 215, 220, 220, 222, 220, 219, 217, 221, 220, 219, 219, 217, 219, 216, 220, 218, 222, 218, 221, 220, 218, 216, 218, 217, 219, 220, 219, 219, 220, 220, 219, 220, 216, 217, 216, 216, 219, 218, 217, 219, 220, 216, 218, 221, 219, 217, 216, 220, 221, 222, 220, 218, 220, 224, 222, 221, 220, 217, 217, 218, 218, 214, 211, 216, 218, 217, 214, 219, 216, 220, 216, 218, 215, 215, 215, 213, 218, 217, 214, 209, 202, 152, 203, 201, 198, 200, 91, 193, 198, 195, 197, 196, 195, 201, 197, 202, 201, 203, 202, 206, 206, 209, 212, 210, 211, 207, 209, 209, 205, 210, 207, 211, 210, 212, 209, 210, 210, 209, 209, 212, 213, 214, 212, 215, 210, 212, 212, 212, 215, 213, 214, 215, 213, 216, 218, 214, 217, 218, 218, 217, 215, 217, 218, 218, 219, 217, 217, 218, 217, 223, 216, 218, 218, 218, 220, 220, 218, 217, 215, 216, 219, 213, 216, 216, 220, 219, 217, 220, 218, 218, 218, 218, 219, 217, 218, 217, 220, 222, 221, 219, 219, 220, 220, 223, 219, 221, 219, 221, 223, 220, 218, 219, 222, 221, 220, 222, 220, 223, 222, 222, 219, 218, 219, 219, 222, 219, 220, 219, 218, 219, 219, 219, 218, 219, 219, 219, 217, 219, 222, 222, 223, 224, 223, 223, 224, 223, 225, 222, 222, 220, 219, 221, 223, 220, 220, 219, 221, 223, 223, 223, 222, 222, 222, 224, 222, 221, 221, 221, 220, 224, 221, 220, 218, 221, 222, 221, 217, 218, 220, 224, 219, 218, 217, 219, 223, 220, 219, 220, 217, 216, 220, 221, 219, 220, 221, 219, 219, 217, 218, 220, 215, 220, 218, 217, 221, 222, 221, 218, 218, 215, 215, 217, 218, 218, 218, 217, 219, 217, 220, 221, 218, 220, 221, 219, 222, 224, 218, 217, 218, 220, 221, 221, 221, 220, 222, 218, 220, 215, 213, 218, 220, 219, 219, 218, 215, 218, 216, 220, 218, 215, 215, 214, 220, 216, 215, 214, 206, 155, 200, 199, 195, 199, 109, 197, 202, 197, 197, 195, 199, 203, 202, 204, 200, 203, 208, 207, 207, 206, 210, 211, 210, 207, 207, 205, 206, 208, 215, 211, 210, 210, 212, 211, 208, 208, 208, 212, 209, 215, 212, 213, 212, 210, 215, 211, 212, 212, 213, 212, 217, 216, 216, 217, 215, 219, 217, 216, 215, 216, 216, 217, 219, 218, 219, 218, 219, 221, 217, 217, 219, 218, 221, 220, 218, 218, 218, 218, 218, 216, 216, 217, 220, 221, 220, 221, 219, 215, 217, 220, 216, 219, 217, 217, 221, 220, 221, 219, 221, 220, 221, 222, 219, 221, 221, 223, 224, 223, 223, 221, 221, 222, 221, 222, 222, 220, 223, 221, 220, 218, 219, 219, 223, 220, 219, 220, 218, 221, 219, 221, 218, 220, 223, 222, 221, 218, 221, 222, 220, 222, 225, 221, 224, 223, 222, 224, 222, 221, 221, 221, 219, 220, 222, 221, 220, 222, 223, 221, 224, 221, 223, 223, 224, 220, 222, 221, 221, 225, 222, 220, 217, 220, 221, 223, 219, 219, 222, 223, 222, 218, 221, 219, 219, 218, 219, 221, 219, 220, 219, 221, 221, 220, 219, 219, 219, 221, 218, 219, 217, 221, 222, 220, 222, 220, 219, 218, 220, 214, 218, 216, 220, 221, 220, 217, 219, 217, 221, 220, 218, 221, 219, 222, 224, 221, 218, 216, 219, 219, 222, 219, 219, 221, 222, 221, 221, 217, 217, 219, 219, 217, 218, 218, 217, 219, 217, 222, 216, 217, 217, 219, 218, 215, 220, 215, 206, 175, 203, 197, 199, 200, 97, 198, 201, 198, 198, 195, 200, 200, 203, 202, 203, 206, 209, 205, 207, 206, 204, 209, 206, 211, 208, 206, 208, 208, 213, 215, 209, 212, 208, 214, 212, 211, 212, 207, 211, 212, 212, 211, 212, 212, 213, 213, 214, 218, 216, 216, 213, 217, 214, 217, 219, 218, 217, 218, 217, 216, 213, 216, 218, 218, 219, 218, 220, 220, 219, 219, 220, 218, 221, 221, 220, 220, 220, 220, 220, 216, 217, 219, 218, 221, 220, 220, 219, 217, 217, 219, 218, 222, 222, 223, 224, 222, 223, 221, 217, 220, 222, 222, 223, 220, 221, 223, 225, 223, 223, 223, 221, 222, 221, 220, 222, 220, 224, 224, 223, 221, 218, 218, 222, 222, 220, 219, 220, 217, 222, 223, 217, 217, 219, 221, 221, 220, 216, 222, 222, 224, 225, 222, 224, 223, 224, 224, 222, 217, 222, 223, 221, 222, 220, 222, 222, 224, 225, 220, 224, 221, 224, 224, 224, 221, 219, 221, 224, 222, 222, 218, 218, 223, 223, 224, 221, 220, 222, 222, 222, 219, 217, 217, 220, 219, 223, 218, 220, 221, 221, 222, 222, 218, 222, 221, 220, 222, 219, 218, 219, 224, 223, 220, 222, 222, 221, 221, 219, 215, 215, 218, 224, 220, 220, 218, 218, 219, 223, 223, 220, 221, 219, 225, 222, 223, 217, 222, 221, 221, 220, 220, 221, 219, 220, 221, 222, 221, 219, 219, 220, 217, 217, 218, 217, 217, 218, 217, 214, 218, 219, 219, 218, 218, 221, 215, 206, 189, 206, 199, 196, 202, 98, 195, 198, 200, 195, 197, 198, 200, 201, 200, 203, 202, 206, 206, 207, 206, 207, 208, 208, 206, 209, 207, 207, 208, 211, 212, 208, 211, 207, 213, 212, 209, 209, 211, 213, 214, 210, 213, 211, 213, 216, 215, 218, 219, 214, 216, 217, 218, 216, 215, 219, 215, 218, 220, 220, 216, 222, 218, 219, 219, 217, 219, 221, 222, 218, 217, 221, 218, 223, 220, 222, 218, 219, 217, 220, 220, 220, 218, 220, 220, 220, 218, 220, 217, 222, 220, 221, 221, 220, 222, 224, 223, 222, 220, 220, 220, 223, 224, 221, 221, 222, 225, 222, 222, 222, 223, 223, 224, 221, 220, 224, 221, 225, 224, 224, 219, 221, 220, 223, 222, 220, 219, 219, 220, 221, 221, 220, 219, 219, 222, 220, 218, 221, 223, 222, 225, 226, 225, 223, 223, 222, 225, 223, 222, 225, 223, 221, 224, 219, 223, 221, 226, 225, 223, 222, 222, 223, 226, 224, 223, 222, 222, 225, 221, 222, 223, 220, 222, 221, 220, 219, 220, 221, 221, 222, 221, 217, 217, 223, 221, 223, 220, 221, 222, 222, 219, 219, 218, 218, 221, 221, 221, 222, 219, 220, 224, 222, 220, 220, 221, 220, 218, 219, 218, 220, 220, 224, 222, 222, 219, 220, 220, 223, 221, 222, 221, 219, 222, 220, 224, 222, 221, 222, 219, 223, 222, 221, 220, 220, 224, 223, 223, 224, 220, 222, 221, 217, 221, 217, 220, 219, 215, 214, 218, 217, 219, 222, 220, 221, 214, 212, 189, 201, 200, 201, 203, 99, 198, 204, 205, 197, 199, 200, 202, 203, 202, 207, 208, 207, 207, 205, 199, 205, 208, 205, 205, 209, 207, 209, 211, 211, 210, 208, 208, 210, 212, 213, 207, 207, 212, 211, 215, 212, 215, 214, 215, 214, 217, 218, 216, 218, 216, 215, 215, 217, 215, 214, 217, 220, 220, 219, 217, 220, 219, 219, 217, 219, 220, 220, 221, 220, 217, 220, 218, 222, 220, 220, 219, 221, 217, 221, 219, 216, 221, 220, 221, 220, 221, 221, 220, 219, 220, 220, 222, 221, 223, 224, 225, 223, 220, 219, 221, 225, 224, 224, 223, 223, 225, 225, 224, 222, 221, 220, 222, 221, 222, 224, 221, 226, 224, 223, 219, 219, 220, 220, 220, 221, 220, 220, 223, 221, 221, 217, 220, 222, 223, 221, 220, 223, 224, 224, 224, 224, 224, 224, 223, 224, 223, 224, 222, 223, 223, 225, 222, 221, 224, 220, 222, 225, 224, 223, 221, 223, 226, 222, 223, 222, 222, 221, 224, 223, 222, 223, 223, 222, 223, 221, 221, 219, 224, 221, 222, 220, 220, 222, 221, 221, 221, 223, 222, 223, 219, 220, 219, 218, 220, 220, 222, 224, 221, 221, 222, 223, 223, 222, 218, 223, 220, 216, 219, 219, 218, 222, 223, 219, 221, 222, 224, 224, 224, 221, 220, 220, 222, 222, 224, 221, 221, 219, 222, 221, 223, 221, 220, 220, 225, 219, 222, 221, 220, 222, 220, 218, 218, 217, 215, 222, 215, 216, 217, 215, 220, 220, 222, 217, 214, 209, 193, 204, 204, 197, 203, 102, 192, 201, 202, 203, 201, 201, 201, 204, 205, 205, 206, 206, 207, 206, 203, 209, 205, 208, 207, 211, 210, 209, 208, 207, 212, 209, 209, 213, 210, 212, 212, 210, 212, 212, 214, 213, 216, 216, 213, 214, 215, 216, 217, 220, 217, 215, 218, 213, 215, 215, 218, 220, 221, 220, 217, 222, 221, 220, 220, 221, 220, 219, 221, 221, 219, 221, 219, 221, 221, 217, 216, 219, 220, 222, 219, 219, 220, 221, 222, 219, 222, 222, 221, 220, 221, 221, 221, 223, 225, 225, 223, 221, 220, 220, 222, 225, 225, 224, 224, 221, 225, 225, 226, 223, 222, 223, 224, 224, 222, 224, 225, 225, 227, 223, 223, 222, 220, 221, 222, 222, 221, 218, 222, 220, 218, 220, 221, 222, 222, 221, 222, 222, 224, 224, 225, 223, 221, 223, 222, 225, 224, 224, 223, 223, 224, 221, 221, 219, 223, 223, 225, 226, 225, 223, 222, 225, 224, 223, 223, 223, 225, 226, 225, 223, 225, 221, 223, 223, 223, 221, 221, 220, 224, 223, 220, 221, 220, 223, 223, 221, 222, 221, 223, 223, 221, 221, 220, 223, 221, 221, 222, 221, 221, 220, 222, 223, 224, 219, 221, 223, 221, 217, 222, 222, 221, 225, 223, 222, 221, 223, 223, 223, 224, 223, 223, 220, 220, 223, 222, 220, 223, 223, 222, 222, 219, 221, 221, 221, 225, 223, 222, 220, 220, 222, 218, 220, 218, 217, 214, 220, 218, 216, 217, 218, 220, 218, 218, 218, 212, 205, 186, 208, 203, 198, 201, 89, 191, 204, 202, 202, 200, 203, 203, 204, 203, 205, 203, 205, 206, 205, 203, 205, 207, 208, 207, 212, 208, 210, 210, 209, 209, 207, 211, 212, 213, 208, 212, 213, 212, 210, 213, 216, 217, 211, 213, 214, 216, 217, 215, 218, 219, 219, 218, 217, 218, 214, 217, 220, 221, 223, 217, 219, 221, 222, 221, 223, 219, 220, 222, 222, 221, 219, 220, 224, 221, 221, 218, 220, 222, 222, 222, 220, 218, 219, 220, 218, 223, 223, 220, 219, 221, 223, 222, 223, 223, 223, 225, 219, 220, 219, 223, 222, 222, 224, 225, 224, 225, 225, 226, 223, 221, 223, 223, 225, 223, 223, 225, 226, 224, 225, 221, 222, 222, 221, 223, 220, 221, 220, 222, 222, 223, 222, 221, 223, 222, 224, 225, 222, 221, 224, 225, 224, 223, 223, 221, 222, 224, 223, 223, 224, 222, 224, 223, 223, 224, 225, 226, 225, 224, 224, 223, 226, 225, 225, 223, 225, 226, 227, 224, 226, 224, 225, 224, 221, 223, 222, 222, 222, 223, 222, 222, 221, 222, 221, 225, 222, 222, 221, 222, 224, 223, 223, 219, 222, 224, 220, 223, 223, 223, 220, 224, 222, 222, 222, 222, 224, 222, 224, 220, 220, 225, 224, 223, 223, 222, 221, 224, 223, 224, 222, 221, 221, 223, 221, 223, 221, 220, 222, 222, 221, 219, 219, 221, 218, 223, 224, 222, 221, 223, 222, 221, 218, 218, 216, 217, 219, 215, 217, 219, 220, 222, 219, 225, 219, 214, 208, 185, 206, 205, 201, 200, 94, 193, 203, 204, 204, 203, 205, 202, 203, 205, 207, 204, 207, 207, 204, 207, 204, 210, 207, 208, 209, 207, 207, 206, 208, 208, 213, 212, 209, 212, 212, 211, 214, 211, 212, 214, 214, 215, 216, 215, 214, 218, 218, 216, 219, 218, 218, 217, 219, 217, 217, 218, 221, 219, 219, 220, 220, 221, 220, 220, 222, 219, 223, 221, 223, 223, 222, 221, 223, 220, 220, 218, 221, 222, 222, 221, 221, 220, 219, 220, 218, 221, 223, 224, 222, 220, 224, 224, 224, 222, 222, 227, 220, 220, 221, 223, 225, 225, 224, 225, 224, 226, 224, 224, 225, 223, 224, 223, 222, 224, 222, 224, 222, 223, 222, 222, 223, 224, 226, 223, 224, 223, 222, 221, 224, 225, 221, 224, 224, 222, 225, 224, 223, 223, 225, 226, 223, 223, 222, 223, 221, 222, 224, 224, 224, 224, 226, 226, 225, 225, 226, 226, 227, 226, 223, 224, 225, 225, 224, 226, 225, 225, 227, 226, 225, 225, 222, 222, 224, 225, 224, 222, 221, 221, 220, 222, 222, 225, 224, 223, 224, 221, 222, 223, 225, 224, 222, 222, 224, 225, 223, 224, 222, 222, 223, 224, 224, 224, 222, 222, 224, 222, 222, 223, 220, 223, 221, 223, 223, 222, 224, 224, 224, 226, 224, 222, 220, 223, 220, 225, 222, 221, 223, 222, 224, 223, 222, 219, 220, 222, 226, 222, 224, 224, 219, 221, 221, 220, 216, 218, 217, 218, 217, 219, 222, 220, 222, 223, 220, 215, 207, 190, 203, 198, 196, 200, 97, 199, 205, 207, 205, 203, 206, 205, 205, 204, 206, 204, 207, 205, 210, 211, 208, 211, 210, 212, 211, 203, 209, 204, 207, 207, 209, 209, 207, 213, 211, 214, 213, 212, 209, 214, 215, 219, 216, 214, 216, 217, 218, 221, 220, 218, 219, 215, 218, 216, 217, 217, 221, 222, 223, 222, 220, 222, 220, 222, 222, 221, 223, 222, 222, 220, 220, 220, 223, 220, 219, 220, 220, 221, 218, 222, 219, 220, 220, 224, 224, 224, 224, 223, 222, 222, 226, 224, 223, 224, 224, 225, 224, 219, 221, 223, 226, 222, 225, 224, 224, 225, 226, 225, 223, 224, 223, 224, 222, 224, 224, 224, 223, 223, 222, 224, 224, 220, 225, 224, 224, 222, 224, 222, 225, 225, 224, 225, 224, 223, 225, 223, 223, 225, 227, 227, 223, 225, 221, 225, 223, 223, 223, 224, 226, 226, 226, 227, 226, 226, 226, 227, 228, 226, 223, 224, 225, 227, 225, 227, 227, 225, 227, 225, 224, 223, 222, 225, 226, 224, 223, 224, 222, 224, 222, 222, 224, 224, 225, 223, 224, 222, 220, 224, 224, 224, 224, 220, 224, 224, 226, 222, 223, 224, 222, 225, 223, 224, 223, 222, 225, 225, 223, 223, 225, 222, 224, 224, 223, 224, 225, 224, 225, 224, 226, 219, 221, 222, 222, 224, 224, 220, 223, 222, 223, 224, 224, 219, 224, 224, 225, 224, 223, 222, 224, 221, 220, 221, 217, 220, 216, 216, 221, 217, 221, 218, 224, 220, 218, 216, 209, 194, 202, 203, 200, 203, 93, 199, 205, 201, 206, 206, 207, 205, 207, 209, 208, 206, 210, 208, 210, 212, 210, 210, 210, 209, 213, 209, 208, 210, 208, 208, 208, 209, 211, 212, 213, 212, 212, 214, 211, 216, 217, 218, 216, 218, 216, 218, 217, 218, 219, 216, 221, 216, 219, 218, 219, 220, 220, 221, 223, 222, 222, 221, 224, 224, 222, 222, 224, 224, 224, 223, 220, 222, 222, 223, 219, 220, 218, 217, 219, 222, 219, 218, 222, 222, 225, 224, 223, 221, 224, 224, 224, 224, 225, 224, 224, 224, 222, 220, 221, 223, 223, 225, 223, 226, 224, 224, 225, 224, 224, 224, 225, 224, 225, 224, 225, 223, 223, 225, 225, 223, 222, 224, 224, 223, 224, 222, 223, 223, 224, 224, 224, 224, 225, 226, 226, 224, 224, 226, 227, 226, 225, 225, 224, 223, 225, 223, 224, 224, 224, 226, 226, 226, 227, 226, 226, 227, 225, 225, 224, 225, 227, 227, 228, 225, 225, 223, 226, 226, 224, 224, 222, 223, 225, 225, 224, 221, 222, 223, 223, 223, 224, 225, 225, 224, 225, 223, 223, 224, 225, 224, 223, 224, 224, 224, 227, 225, 223, 224, 223, 224, 225, 223, 224, 224, 223, 225, 223, 222, 221, 223, 222, 222, 222, 223, 223, 222, 226, 224, 224, 221, 222, 222, 223, 226, 221, 222, 223, 224, 224, 223, 222, 217, 219, 223, 224, 225, 223, 224, 222, 223, 219, 219, 220, 217, 219, 215, 217, 215, 220, 220, 223, 220, 220, 218, 210, 193, 203, 203, 201, 202, 100, 198, 207, 202, 202, 206, 207, 204, 207, 211, 207, 210, 211, 211, 210, 212, 213, 209, 212, 211, 212, 212, 210, 210, 212, 210, 209, 210, 210, 212, 210, 215, 213, 213, 217, 217, 218, 217, 215, 218, 217, 218, 223, 220, 217, 216, 220, 215, 220, 220, 220, 222, 222, 220, 221, 221, 218, 223, 223, 223, 223, 224, 223, 222, 223, 222, 221, 222, 221, 222, 217, 220, 220, 219, 222, 222, 218, 219, 222, 224, 224, 223, 220, 224, 222, 225, 225, 225, 224, 223, 225, 223, 225, 220, 221, 224, 225, 224, 224, 225, 223, 225, 224, 227, 224, 224, 226, 227, 227, 225, 224, 224, 221, 224, 225, 224, 222, 224, 225, 226, 224, 224, 225, 222, 225, 225, 224, 223, 224, 225, 226, 224, 225, 227, 229, 228, 229, 225, 224, 223, 222, 224, 223, 223, 223, 224, 225, 227, 227, 225, 226, 226, 229, 227, 226, 224, 226, 224, 225, 226, 225, 227, 228, 228, 225, 224, 224, 225, 224, 224, 225, 223, 224, 226, 224, 225, 225, 224, 225, 226, 227, 223, 222, 225, 225, 224, 224, 222, 222, 223, 226, 224, 222, 223, 224, 223, 225, 226, 224, 224, 224, 223, 224, 220, 220, 219, 224, 223, 224, 224, 225, 224, 224, 223, 224, 223, 221, 222, 218, 224, 220, 223, 223, 223, 224, 225, 222, 220, 221, 224, 224, 225, 224, 223, 224, 222, 222, 219, 217, 219, 220, 216, 222, 220, 221, 220, 219, 222, 219, 214, 208, 193, 204, 203, 204, 204, 102, 200, 203, 202, 203, 207, 209, 207, 210, 208, 211, 208, 208, 210, 210, 211, 215, 208, 215, 213, 216, 212, 209, 212, 210, 211, 210, 210, 210, 214, 212, 215, 211, 213, 218, 216, 219, 218, 218, 216, 216, 220, 221, 220, 217, 218, 216, 217, 215, 221, 218, 222, 220, 225, 224, 221, 222, 224, 223, 223, 221, 223, 223, 222, 223, 221, 220, 219, 221, 222, 217, 219, 219, 220, 222, 219, 221, 221, 220, 221, 223, 225, 223, 224, 225, 228, 225, 225, 224, 225, 227, 225, 226, 222, 223, 224, 226, 223, 225, 227, 227, 225, 226, 226, 222, 224, 227, 226, 226, 226, 223, 223, 223, 224, 225, 224, 224, 224, 223, 226, 224, 225, 224, 225, 224, 227, 222, 223, 224, 224, 225, 225, 226, 225, 228, 228, 228, 227, 226, 224, 227, 224, 226, 225, 226, 225, 227, 228, 227, 225, 226, 229, 228, 227, 224, 225, 227, 224, 227, 226, 227, 226, 227, 229, 226, 224, 226, 222, 226, 226, 223, 223, 224, 225, 224, 227, 225, 223, 227, 226, 227, 223, 222, 223, 224, 225, 223, 224, 222, 223, 226, 226, 224, 225, 223, 225, 224, 225, 224, 223, 226, 225, 224, 221, 223, 220, 224, 224, 227, 224, 223, 224, 224, 224, 222, 225, 223, 225, 226, 223, 222, 224, 225, 223, 223, 224, 222, 220, 224, 225, 224, 225, 223, 223, 224, 222, 222, 220, 220, 219, 220, 221, 219, 223, 221, 222, 221, 222, 217, 217, 208, 194, 205, 201, 202, 203, 102, 198, 205, 202, 201, 206, 206, 208, 212, 208, 210, 205, 206, 210, 211, 214, 213, 213, 214, 211, 212, 213, 211, 210, 213, 214, 211, 214, 212, 212, 213, 212, 214, 215, 219, 217, 218, 219, 217, 217, 219, 219, 219, 219, 220, 219, 220, 220, 218, 219, 218, 222, 222, 223, 223, 222, 224, 221, 224, 221, 222, 224, 221, 224, 223, 221, 221, 220, 220, 220, 218, 219, 220, 222, 221, 219, 222, 222, 222, 222, 225, 224, 224, 223, 224, 225, 224, 225, 226, 224, 226, 225, 224, 225, 225, 226, 226, 226, 226, 227, 226, 225, 226, 226, 224, 224, 224, 226, 225, 224, 225, 223, 226, 226, 226, 224, 224, 226, 226, 226, 226, 223, 224, 226, 224, 225, 224, 224, 225, 224, 226, 225, 225, 226, 228, 229, 229, 225, 227, 226, 226, 226, 227, 227, 225, 226, 228, 226, 226, 224, 225, 229, 227, 226, 221, 223, 225, 225, 226, 227, 227, 226, 228, 227, 228, 225, 227, 226, 226, 224, 223, 225, 223, 224, 224, 224, 226, 224, 226, 226, 225, 225, 224, 223, 224, 225, 224, 224, 224, 224, 227, 227, 224, 223, 221, 226, 226, 225, 223, 223, 225, 225, 224, 225, 222, 223, 223, 225, 225, 223, 224, 224, 224, 223, 224, 225, 223, 224, 224, 223, 223, 225, 227, 222, 224, 224, 225, 223, 224, 225, 226, 224, 225, 220, 225, 224, 222, 219, 219, 219, 220, 222, 221, 223, 222, 222, 221, 222, 220, 213, 208, 195, 207, 200, 201, 202, 99, 197, 203, 202, 204, 206, 204, 207, 211, 214, 212, 209, 206, 207, 213, 213, 215, 214, 215, 216, 212, 214, 215, 214, 213, 214, 211, 212, 213, 214, 216, 213, 213, 216, 217, 219, 220, 216, 218, 216, 218, 218, 221, 220, 221, 220, 221, 221, 220, 221, 222, 223, 223, 224, 222, 220, 224, 224, 224, 222, 223, 223, 221, 224, 223, 223, 223, 221, 223, 220, 220, 219, 219, 222, 223, 222, 223, 220, 221, 226, 224, 224, 224, 223, 226, 227, 226, 226, 226, 226, 227, 227, 224, 226, 225, 227, 226, 226, 226, 228, 226, 226, 227, 225, 226, 224, 224, 226, 225, 224, 224, 225, 226, 227, 227, 225, 224, 226, 224, 225, 225, 225, 225, 225, 225, 225, 225, 226, 226, 224, 224, 227, 225, 228, 229, 229, 228, 227, 227, 228, 226, 227, 227, 225, 225, 225, 226, 224, 225, 224, 225, 228, 229, 227, 224, 222, 226, 223, 227, 225, 225, 227, 227, 228, 228, 226, 226, 226, 227, 225, 221, 225, 222, 222, 225, 224, 224, 224, 225, 226, 227, 225, 224, 224, 223, 224, 224, 223, 224, 222, 226, 226, 226, 221, 221, 227, 226, 224, 224, 223, 225, 224, 227, 224, 219, 224, 226, 225, 225, 222, 222, 225, 223, 222, 225, 224, 225, 222, 224, 216, 220, 223, 223, 222, 226, 225, 224, 222, 225, 224, 224, 220, 221, 221, 224, 224, 221, 224, 221, 222, 221, 222, 221, 221, 219, 223, 220, 219, 217, 212, 205, 195, 207, 204, 202, 201, 105, 198, 204, 202, 203, 205, 207, 209, 210, 213, 211, 205, 208, 212, 212, 211, 215, 216, 213, 214, 211, 212, 213, 215, 214, 214, 211, 213, 213, 216, 215, 216, 215, 217, 217, 218, 220, 220, 220, 220, 220, 219, 219, 221, 222, 220, 221, 223, 221, 219, 223, 224, 222, 221, 223, 221, 221, 224, 222, 223, 224, 223, 223, 226, 225, 223, 223, 224, 224, 224, 219, 221, 219, 222, 223, 224, 222, 223, 222, 226, 226, 226, 223, 225, 226, 226, 227, 225, 225, 225, 227, 226, 223, 225, 224, 226, 225, 224, 225, 227, 226, 227, 227, 225, 225, 226, 227, 226, 226, 224, 225, 226, 226, 226, 226, 225, 223, 225, 227, 225, 226, 224, 226, 227, 226, 227, 226, 227, 227, 228, 226, 226, 227, 226, 228, 229, 229, 228, 226, 228, 227, 229, 228, 226, 224, 226, 227, 227, 227, 228, 228, 228, 228, 227, 226, 224, 225, 226, 226, 227, 225, 227, 227, 228, 229, 227, 226, 225, 227, 225, 224, 222, 222, 225, 224, 225, 224, 224, 227, 227, 226, 225, 224, 224, 225, 226, 223, 223, 224, 225, 228, 227, 225, 223, 224, 225, 226, 223, 222, 224, 223, 226, 226, 223, 224, 222, 223, 226, 224, 223, 223, 224, 225, 225, 224, 224, 224, 225, 227, 221, 219, 225, 224, 225, 225, 225, 224, 224, 227, 225, 224, 220, 223, 222, 222, 225, 223, 219, 222, 220, 222, 222, 220, 220, 223, 222, 221, 222, 220, 214, 205, 198, 203, 207, 201, 205, 92, 196, 203, 205, 204, 204, 212, 212, 211, 213, 208, 203, 207, 212, 213, 214, 216, 216, 213, 212, 214, 214, 213, 216, 214, 214, 213, 212, 213, 217, 214, 216, 214, 218, 219, 217, 219, 220, 222, 220, 219, 218, 220, 220, 223, 219, 222, 221, 220, 221, 222, 224, 224, 224, 221, 222, 222, 222, 222, 223, 223, 222, 224, 226, 225, 225, 224, 225, 224, 224, 222, 218, 221, 224, 223, 223, 225, 222, 225, 226, 227, 226, 224, 225, 226, 226, 226, 226, 225, 227, 227, 225, 226, 225, 226, 225, 224, 227, 226, 227, 226, 226, 227, 227, 225, 226, 227, 225, 225, 226, 226, 226, 227, 227, 227, 225, 224, 224, 228, 225, 226, 226, 225, 226, 227, 227, 225, 228, 228, 228, 226, 227, 227, 226, 227, 228, 227, 228, 228, 228, 228, 228, 226, 227, 224, 229, 227, 227, 225, 226, 227, 227, 230, 228, 226, 226, 226, 224, 227, 226, 224, 226, 226, 229, 228, 227, 227, 226, 225, 227, 223, 223, 223, 225, 226, 226, 226, 226, 227, 227, 225, 226, 225, 224, 226, 225, 223, 224, 223, 225, 225, 227, 223, 224, 225, 225, 225, 227, 224, 224, 222, 227, 225, 225, 225, 225, 226, 225, 225, 224, 222, 223, 225, 224, 225, 225, 225, 227, 227, 221, 223, 224, 227, 227, 226, 225, 225, 224, 225, 225, 225, 223, 222, 221, 224, 225, 223, 220, 220, 223, 220, 221, 221, 220, 224, 221, 224, 220, 218, 213, 207, 199, 204, 202, 203, 209, 120, 201, 206, 204, 205, 205, 209, 211, 212, 212, 210, 206, 208, 209, 214, 215, 212, 212, 211, 211, 215, 214, 216, 215, 214, 214, 214, 213, 216, 218, 215, 213, 216, 218, 219, 222, 218, 222, 220, 222, 221, 221, 219, 222, 224, 219, 223, 222, 221, 219, 221, 221, 226, 224, 223, 220, 222, 221, 223, 222, 224, 221, 223, 225, 225, 225, 224, 224, 225, 224, 223, 223, 221, 224, 223, 222, 222, 222, 225, 225, 226, 226, 224, 223, 225, 227, 225, 224, 224, 226, 227, 226, 226, 223, 227, 227, 226, 227, 227, 226, 226, 227, 226, 226, 224, 225, 226, 225, 226, 224, 225, 224, 225, 226, 227, 226, 226, 227, 227, 225, 226, 225, 225, 226, 229, 227, 226, 227, 226, 227, 226, 226, 226, 227, 226, 230, 229, 227, 228, 228, 229, 229, 227, 226, 225, 227, 226, 228, 226, 225, 229, 229, 227, 228, 226, 226, 229, 227, 227, 225, 227, 227, 228, 229, 228, 228, 228, 228, 226, 227, 224, 221, 223, 225, 225, 225, 226, 227, 228, 226, 227, 227, 225, 224, 227, 226, 225, 223, 223, 223, 226, 226, 226, 222, 225, 227, 224, 227, 225, 224, 224, 226, 226, 224, 226, 224, 228, 225, 222, 221, 222, 221, 226, 226, 224, 225, 227, 226, 227, 225, 225, 223, 226, 227, 225, 226, 223, 224, 226, 226, 225, 224, 224, 224, 224, 224, 223, 222, 222, 220, 219, 220, 223, 221, 222, 222, 222, 220, 220, 217, 208, 201, 204, 204, 202, 208, 124, 208, 201, 204, 210, 207, 211, 207, 215, 215, 214, 210, 208, 210, 212, 213, 211, 212, 212, 209, 216, 214, 214, 212, 214, 216, 214, 211, 216, 215, 212, 216, 218, 218, 218, 221, 221, 219, 220, 221, 222, 222, 219, 221, 224, 221, 224, 222, 224, 221, 221, 222, 224, 221, 221, 222, 219, 222, 223, 224, 224, 221, 223, 224, 224, 225, 224, 224, 222, 222, 223, 224, 221, 223, 222, 225, 223, 225, 225, 226, 225, 226, 225, 224, 227, 226, 224, 223, 225, 226, 226, 227, 227, 226, 227, 226, 227, 227, 227, 226, 227, 227, 227, 228, 226, 225, 227, 227, 227, 225, 225, 222, 226, 227, 227, 225, 226, 227, 226, 227, 226, 224, 225, 227, 227, 227, 224, 226, 226, 225, 227, 227, 227, 226, 228, 227, 228, 228, 227, 228, 229, 228, 228, 227, 225, 227, 228, 225, 226, 226, 227, 229, 227, 228, 228, 228, 228, 227, 228, 227, 226, 228, 227, 227, 228, 228, 227, 225, 225, 228, 225, 223, 224, 225, 224, 225, 225, 226, 226, 225, 224, 226, 225, 222, 226, 227, 225, 224, 220, 223, 223, 224, 227, 225, 226, 225, 225, 223, 223, 222, 225, 224, 225, 226, 226, 225, 225, 224, 221, 223, 222, 223, 226, 227, 224, 224, 226, 226, 227, 226, 226, 224, 228, 227, 227, 227, 225, 224, 226, 226, 227, 226, 225, 227, 225, 226, 221, 220, 220, 223, 222, 220, 221, 221, 221, 222, 222, 223, 219, 217, 209, 204, 207, 205, 202, 209, 135, 204, 203, 207, 208, 212, 210, 212, 214, 215, 213, 209, 209, 212, 212, 213, 212, 210, 211, 210, 213, 213, 213, 215, 215, 216, 213, 214, 213, 217, 214, 217, 217, 215, 216, 222, 222, 221, 220, 219, 223, 221, 221, 223, 223, 224, 224, 224, 223, 221, 221, 223, 225, 219, 224, 223, 222, 225, 222, 222, 223, 222, 224, 225, 225, 225, 225, 223, 226, 223, 222, 223, 224, 224, 226, 225, 223, 224, 225, 227, 225, 226, 225, 225, 225, 226, 225, 221, 225, 225, 224, 227, 225, 227, 227, 227, 227, 228, 227, 226, 225, 227, 227, 228, 227, 225, 226, 227, 227, 223, 225, 223, 226, 227, 226, 225, 226, 227, 225, 227, 226, 226, 226, 228, 228, 228, 226, 226, 226, 228, 226, 226, 227, 227, 229, 228, 228, 228, 227, 227, 228, 229, 228, 227, 227, 229, 227, 223, 225, 226, 227, 226, 229, 228, 227, 227, 227, 227, 228, 226, 228, 228, 228, 228, 228, 228, 227, 226, 228, 227, 225, 225, 222, 224, 224, 227, 225, 226, 226, 226, 227, 223, 225, 226, 225, 226, 226, 224, 224, 224, 222, 226, 227, 226, 226, 224, 225, 225, 223, 224, 224, 223, 224, 223, 224, 224, 226, 226, 224, 225, 223, 225, 225, 227, 225, 225, 226, 225, 228, 227, 225, 226, 227, 228, 228, 227, 225, 224, 226, 224, 225, 225, 225, 228, 226, 226, 224, 223, 222, 221, 222, 224, 221, 222, 222, 221, 222, 219, 217, 214, 211, 206, 208, 200, 204, 210, 120, 202, 207, 208, 208, 210, 208, 210, 209, 212, 212, 211, 211, 212, 214, 213, 208, 211, 214, 213, 213, 211, 213, 215, 210, 212, 215, 217, 214, 218, 217, 221, 218, 217, 218, 225, 221, 222, 222, 219, 223, 223, 224, 224, 225, 225, 225, 226, 224, 224, 223, 225, 225, 221, 224, 223, 224, 224, 226, 224, 224, 222, 224, 224, 224, 226, 226, 223, 224, 224, 224, 224, 225, 226, 225, 226, 225, 224, 225, 225, 225, 225, 224, 225, 226, 226, 225, 225, 224, 225, 225, 224, 226, 226, 225, 226, 227, 228, 225, 226, 227, 227, 227, 228, 227, 226, 228, 229, 227, 226, 225, 225, 228, 226, 226, 226, 227, 228, 225, 226, 227, 226, 227, 227, 228, 228, 228, 228, 228, 230, 226, 227, 227, 228, 228, 228, 228, 228, 228, 227, 228, 228, 228, 228, 228, 228, 228, 225, 224, 225, 225, 228, 229, 228, 228, 228, 228, 230, 230, 228, 227, 226, 227, 229, 229, 225, 227, 228, 224, 226, 227, 223, 225, 226, 225, 225, 224, 224, 224, 226, 227, 224, 225, 224, 225, 227, 227, 225, 223, 222, 224, 225, 225, 223, 224, 225, 226, 225, 224, 223, 224, 226, 225, 222, 224, 225, 227, 228, 226, 224, 224, 224, 227, 226, 225, 225, 227, 224, 228, 226, 225, 227, 226, 228, 227, 226, 224, 226, 225, 226, 225, 225, 225, 225, 224, 227, 225, 223, 223, 219, 221, 221, 222, 221, 223, 220, 218, 218, 215, 219, 212, 205, 207, 202, 201, 206, 112, 204, 205, 211, 207, 211, 208, 210, 208, 211, 212, 213, 212, 211, 214, 214, 212, 213, 215, 210, 212, 211, 212, 212, 213, 217, 215, 216, 213, 217, 220, 220, 219, 215, 217, 223, 224, 221, 222, 222, 224, 226, 224, 224, 224, 225, 223, 227, 225, 223, 224, 226, 224, 223, 222, 224, 227, 225, 226, 225, 224, 224, 226, 225, 223, 227, 224, 224, 224, 224, 222, 224, 224, 224, 225, 227, 225, 226, 227, 228, 226, 225, 225, 225, 226, 226, 225, 226, 224, 225, 226, 226, 226, 228, 226, 228, 227, 229, 227, 226, 227, 227, 227, 227, 227, 226, 225, 229, 227, 226, 227, 226, 229, 227, 227, 226, 228, 227, 229, 226, 226, 227, 226, 228, 227, 228, 227, 228, 228, 230, 228, 228, 225, 227, 228, 229, 229, 229, 228, 228, 228, 227, 229, 228, 228, 229, 228, 227, 226, 225, 228, 229, 229, 228, 228, 227, 228, 230, 229, 229, 225, 226, 225, 228, 228, 225, 226, 227, 226, 225, 226, 225, 224, 226, 227, 225, 223, 225, 226, 224, 225, 221, 224, 225, 224, 226, 223, 224, 223, 225, 226, 225, 225, 224, 225, 226, 226, 225, 222, 224, 223, 226, 224, 225, 225, 225, 227, 228, 227, 226, 224, 227, 227, 227, 226, 225, 226, 226, 226, 227, 225, 228, 227, 226, 226, 226, 226, 223, 224, 226, 225, 224, 225, 226, 225, 225, 220, 222, 221, 222, 220, 221, 222, 221, 221, 220, 220, 221, 219, 217, 211, 205, 209, 203, 204, 206, 113, 202, 211, 209, 210, 207, 207, 209, 208, 215, 214, 214, 212, 213, 215, 212, 213, 214, 216, 212, 212, 216, 215, 213, 216, 220, 215, 217, 216, 218, 222, 219, 220, 216, 217, 224, 222, 220, 220, 221, 225, 226, 223, 223, 224, 224, 225, 224, 225, 224, 225, 224, 226, 225, 225, 226, 225, 226, 225, 225, 223, 225, 226, 226, 226, 227, 224, 225, 226, 226, 224, 226, 226, 224, 225, 226, 224, 226, 226, 227, 227, 225, 226, 226, 226, 227, 226, 224, 224, 225, 228, 229, 226, 227, 226, 228, 227, 227, 227, 226, 228, 227, 228, 228, 227, 227, 226, 229, 227, 227, 227, 226, 228, 230, 228, 226, 227, 227, 227, 227, 226, 227, 228, 227, 227, 229, 227, 228, 228, 230, 229, 228, 227, 227, 228, 228, 228, 227, 227, 227, 228, 227, 230, 228, 228, 229, 228, 229, 227, 226, 227, 229, 229, 227, 228, 228, 228, 230, 229, 227, 227, 225, 225, 227, 226, 222, 225, 226, 226, 226, 226, 224, 223, 225, 226, 227, 224, 225, 225, 224, 221, 221, 222, 225, 225, 224, 225, 224, 226, 224, 226, 226, 226, 226, 226, 227, 227, 228, 225, 225, 226, 228, 227, 226, 227, 224, 227, 227, 226, 223, 226, 226, 226, 226, 224, 225, 225, 227, 227, 229, 228, 227, 226, 228, 227, 225, 225, 224, 225, 226, 225, 225, 225, 227, 226, 223, 223, 225, 220, 222, 222, 223, 222, 222, 221, 220, 222, 219, 219, 218, 209, 205, 206, 202, 201, 204, 109, 204, 208, 213, 210, 203, 206, 212, 208, 214, 214, 211, 212, 214, 215, 213, 216, 215, 213, 214, 213, 217, 216, 218, 216, 220, 216, 217, 218, 220, 224, 221, 219, 214, 218, 222, 220, 222, 219, 221, 223, 225, 222, 221, 224, 224, 224, 225, 227, 226, 224, 225, 226, 225, 225, 224, 225, 225, 225, 225, 225, 226, 226, 228, 227, 225, 225, 225, 225, 226, 225, 226, 225, 226, 226, 227, 224, 226, 226, 227, 228, 226, 226, 224, 225, 225, 225, 225, 224, 225, 227, 227, 225, 227, 227, 226, 228, 229, 227, 227, 227, 227, 229, 227, 227, 227, 227, 228, 229, 228, 228, 228, 229, 229, 227, 226, 228, 227, 229, 228, 227, 228, 228, 229, 228, 228, 228, 227, 229, 229, 230, 229, 226, 227, 229, 229, 228, 227, 228, 228, 229, 229, 228, 227, 227, 229, 229, 228, 228, 227, 228, 230, 229, 228, 226, 226, 229, 230, 227, 226, 226, 226, 226, 227, 226, 223, 225, 227, 227, 225, 226, 224, 221, 224, 225, 228, 225, 226, 225, 224, 222, 222, 220, 225, 223, 224, 223, 222, 226, 225, 227, 227, 228, 226, 225, 228, 226, 226, 227, 226, 226, 227, 228, 226, 225, 226, 228, 227, 224, 223, 227, 227, 226, 225, 223, 224, 225, 227, 228, 230, 228, 227, 228, 228, 227, 228, 225, 224, 226, 225, 226, 226, 225, 223, 224, 225, 222, 224, 221, 224, 222, 224, 222, 222, 224, 221, 219, 219, 220, 218, 210, 211, 209, 206, 201, 205, 101, 204, 209, 211, 210, 204, 207, 210, 208, 211, 214, 211, 210, 216, 215, 213, 216, 216, 217, 215, 217, 217, 216, 216, 217, 221, 219, 217, 217, 220, 222, 220, 218, 214, 215, 222, 218, 220, 221, 221, 220, 223, 222, 224, 225, 224, 225, 226, 225, 226, 224, 227, 225, 225, 223, 224, 224, 225, 223, 225, 224, 226, 226, 227, 226, 225, 225, 225, 224, 226, 225, 226, 225, 226, 227, 226, 225, 226, 225, 228, 227, 227, 224, 225, 224, 224, 224, 225, 226, 226, 228, 228, 227, 227, 226, 227, 227, 227, 228, 225, 226, 227, 228, 228, 228, 227, 228, 229, 228, 228, 228, 227, 227, 229, 228, 227, 227, 227, 227, 228, 228, 227, 228, 228, 228, 228, 227, 229, 230, 230, 229, 227, 228, 227, 228, 227, 228, 229, 229, 229, 230, 228, 228, 228, 227, 229, 228, 229, 227, 228, 228, 229, 230, 228, 226, 226, 229, 228, 229, 226, 226, 225, 227, 227, 227, 224, 225, 225, 227, 227, 228, 225, 224, 223, 226, 226, 227, 226, 226, 225, 223, 222, 222, 223, 223, 221, 224, 222, 223, 224, 227, 227, 227, 227, 227, 227, 229, 227, 225, 226, 225, 227, 225, 224, 226, 226, 227, 228, 227, 225, 226, 226, 226, 226, 225, 225, 226, 228, 228, 228, 227, 227, 228, 227, 228, 228, 228, 227, 227, 226, 226, 224, 225, 225, 224, 222, 223, 222, 224, 226, 224, 222, 224, 222, 226, 223, 222, 220, 221, 217, 209, 208, 207, 202, 199, 206, 96, 203, 213, 211, 209, 206, 208, 209, 214, 214, 211, 215, 215, 213, 213, 210, 218, 218, 217, 218, 215, 216, 215, 217, 218, 221, 220, 218, 220, 223, 221, 218, 216, 216, 215, 218, 220, 221, 220, 222, 221, 223, 221, 224, 223, 224, 226, 227, 225, 227, 225, 225, 226, 227, 225, 226, 224, 223, 225, 225, 226, 225, 226, 225, 225, 227, 224, 223, 224, 226, 227, 227, 226, 226, 227, 228, 225, 226, 226, 227, 227, 227, 226, 226, 226, 225, 225, 226, 225, 227, 228, 227, 228, 226, 227, 228, 228, 229, 228, 227, 227, 228, 229, 228, 228, 226, 227, 228, 229, 228, 228, 228, 229, 229, 227, 227, 227, 227, 229, 227, 228, 226, 228, 228, 229, 229, 229, 229, 229, 230, 230, 228, 226, 228, 227, 228, 228, 228, 229, 228, 230, 230, 229, 228, 229, 230, 229, 230, 229, 229, 229, 229, 228, 228, 227, 227, 229, 229, 228, 227, 225, 226, 228, 229, 225, 226, 225, 227, 228, 228, 226, 224, 224, 225, 226, 227, 228, 228, 226, 226, 224, 223, 224, 223, 220, 223, 221, 221, 221, 225, 227, 227, 226, 227, 226, 229, 228, 228, 226, 226, 227, 229, 226, 227, 225, 225, 227, 227, 226, 224, 226, 227, 226, 227, 226, 225, 226, 229, 230, 228, 228, 227, 227, 229, 228, 227, 226, 226, 228, 227, 224, 225, 225, 224, 224, 226, 224, 224, 224, 226, 227, 225, 224, 224, 224, 223, 221, 218, 220, 218, 212, 209, 210, 204, 202, 205, 107, 204, 211, 213, 213, 208, 210, 211, 214, 212, 213, 213, 214, 216, 213, 215, 214, 217, 216, 214, 212, 213, 216, 214, 215, 220, 222, 221, 218, 224, 223, 219, 216, 216, 217, 218, 218, 220, 219, 221, 221, 222, 222, 222, 224, 226, 226, 226, 225, 227, 225, 227, 225, 226, 225, 227, 223, 224, 225, 225, 227, 227, 226, 224, 225, 225, 225, 222, 224, 226, 226, 226, 225, 226, 227, 227, 227, 226, 226, 228, 226, 228, 225, 225, 226, 226, 226, 226, 225, 226, 227, 226, 227, 227, 226, 226, 228, 228, 227, 227, 228, 229, 229, 229, 227, 228, 228, 228, 228, 228, 228, 228, 229, 229, 226, 227, 227, 228, 229, 228, 227, 227, 229, 229, 230, 229, 228, 228, 228, 229, 229, 228, 227, 227, 228, 229, 227, 228, 228, 228, 229, 229, 229, 228, 229, 230, 230, 230, 228, 228, 229, 229, 228, 228, 228, 229, 229, 230, 227, 226, 226, 226, 227, 228, 225, 227, 227, 228, 228, 228, 226, 223, 224, 226, 226, 226, 227, 227, 225, 225, 226, 223, 223, 225, 224, 223, 222, 221, 221, 225, 225, 228, 226, 227, 227, 229, 228, 228, 226, 226, 227, 227, 225, 224, 225, 223, 227, 228, 227, 226, 224, 227, 227, 227, 228, 228, 227, 229, 228, 229, 227, 227, 227, 228, 229, 226, 223, 225, 225, 226, 225, 226, 223, 225, 226, 227, 225, 223, 224, 224, 226, 223, 226, 225, 224, 221, 222, 220, 219, 217, 215, 212, 211, 203, 207, 208, 114, 202, 211, 210, 211, 209, 207, 211, 215, 217, 215, 217, 218, 218, 216, 215, 214, 218, 219, 214, 216, 210, 212, 214, 216, 218, 220, 220, 218, 223, 221, 220, 222, 220, 220, 222, 222, 223, 221, 219, 221, 221, 223, 221, 224, 226, 226, 227, 225, 226, 226, 225, 225, 225, 225, 226, 225, 224, 226, 227, 227, 225, 226, 224, 226, 224, 223, 224, 225, 225, 225, 225, 224, 226, 226, 227, 227, 227, 228, 228, 227, 226, 225, 225, 225, 225, 225, 225, 226, 227, 228, 228, 227, 227, 225, 225, 227, 227, 227, 226, 227, 228, 228, 228, 227, 227, 229, 228, 228, 226, 228, 228, 228, 230, 228, 227, 228, 228, 229, 229, 228, 228, 227, 230, 230, 229, 228, 228, 229, 228, 228, 227, 226, 227, 229, 228, 228, 229, 228, 229, 229, 230, 228, 229, 229, 229, 229, 230, 228, 227, 227, 229, 229, 229, 228, 230, 230, 231, 229, 227, 226, 225, 227, 229, 226, 227, 227, 228, 227, 226, 225, 224, 225, 226, 228, 228, 226, 226, 227, 227, 227, 222, 224, 225, 226, 227, 223, 223, 223, 225, 223, 227, 227, 227, 227, 228, 227, 229, 226, 226, 227, 227, 227, 226, 226, 226, 228, 228, 227, 226, 227, 228, 229, 228, 227, 227, 226, 228, 228, 229, 227, 227, 225, 227, 228, 227, 225, 226, 228, 227, 226, 225, 221, 225, 226, 227, 226, 224, 222, 225, 225, 226, 227, 225, 224, 222, 220, 220, 221, 218, 212, 212, 212, 208, 210, 210, 125, 204, 213, 210, 211, 211, 210, 209, 214, 216, 215, 215, 214, 217, 218, 215, 218, 217, 217, 216, 216, 214, 216, 214, 218, 220, 222, 218, 220, 222, 221, 219, 221, 220, 221, 221, 222, 222, 219, 221, 222, 223, 224, 222, 224, 225, 226, 228, 225, 226, 226, 228, 226, 227, 226, 226, 224, 225, 227, 227, 225, 225, 226, 226, 225, 223, 223, 225, 224, 225, 225, 226, 226, 226, 227, 227, 227, 227, 228, 228, 227, 228, 227, 226, 227, 227, 228, 226, 227, 227, 228, 228, 228, 228, 226, 226, 226, 227, 227, 225, 227, 226, 228, 228, 228, 227, 229, 228, 228, 225, 227, 227, 229, 230, 229, 228, 226, 228, 229, 229, 228, 228, 228, 230, 229, 230, 228, 229, 228, 230, 228, 228, 228, 228, 230, 230, 230, 229, 228, 229, 231, 229, 229, 229, 230, 228, 230, 230, 229, 227, 227, 229, 228, 229, 230, 230, 230, 231, 229, 227, 227, 226, 227, 229, 226, 222, 218, 212, 207, 203, 199, 200, 205, 212, 218, 221, 223, 226, 226, 224, 226, 221, 225, 225, 225, 227, 226, 224, 224, 225, 223, 224, 226, 226, 225, 227, 228, 228, 226, 225, 229, 228, 229, 227, 227, 225, 228, 228, 228, 227, 228, 226, 227, 227, 228, 228, 227, 228, 230, 228, 227, 226, 226, 228, 227, 227, 225, 227, 228, 227, 227, 225, 222, 226, 226, 227, 226, 225, 225, 225, 227, 228, 226, 227, 222, 222, 223, 223, 221, 218, 214, 215, 211, 210, 209, 212, 117, 204, 213, 211, 210, 210, 209, 210, 214, 215, 211, 214, 215, 218, 217, 215, 217, 217, 221, 219, 219, 214, 217, 217, 218, 218, 219, 220, 221, 221, 220, 220, 222, 221, 222, 223, 223, 222, 223, 222, 225, 225, 226, 225, 224, 224, 228, 228, 227, 227, 227, 228, 225, 226, 225, 226, 226, 226, 227, 228, 225, 226, 227, 227, 223, 221, 224, 226, 225, 225, 226, 226, 226, 227, 228, 228, 227, 227, 227, 228, 228, 228, 227, 228, 228, 228, 228, 226, 229, 227, 228, 227, 229, 228, 227, 227, 227, 226, 227, 226, 228, 227, 230, 228, 227, 227, 228, 229, 228, 226, 226, 228, 229, 229, 229, 229, 227, 228, 228, 230, 229, 229, 228, 230, 228, 230, 230, 228, 229, 231, 229, 228, 227, 229, 230, 230, 229, 229, 228, 229, 230, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 233, 233, 232, 234, 235, 233, 232, 230, 224, 209, 191, 162, 134, 108, 90, 76, 74, 68, 69, 71, 84, 96, 123, 147, 175, 192, 202, 211, 216, 220, 225, 226, 227, 228, 225, 227, 226, 224, 225, 225, 228, 229, 228, 227, 228, 227, 225, 226, 228, 229, 226, 226, 227, 226, 229, 229, 226, 228, 228, 229, 229, 229, 228, 228, 228, 229, 229, 226, 225, 227, 227, 226, 228, 227, 226, 228, 228, 228, 225, 225, 226, 225, 227, 227, 225, 224, 227, 226, 227, 226, 224, 219, 222, 222, 223, 223, 217, 213, 211, 213, 212, 210, 212, 124, 208, 214, 211, 210, 208, 211, 210, 210, 216, 212, 216, 212, 218, 216, 217, 217, 218, 219, 219, 219, 216, 214, 219, 216, 220, 220, 219, 222, 223, 220, 222, 221, 221, 221, 222, 224, 224, 221, 223, 221, 226, 227, 224, 224, 224, 226, 226, 226, 226, 226, 227, 224, 225, 226, 226, 226, 227, 226, 227, 226, 226, 226, 227, 226, 223, 224, 226, 225, 225, 225, 226, 225, 227, 228, 228, 226, 226, 227, 226, 228, 228, 228, 227, 227, 228, 227, 228, 228, 227, 228, 228, 229, 228, 227, 227, 228, 228, 226, 228, 227, 229, 230, 230, 228, 228, 228, 229, 226, 227, 227, 228, 229, 230, 230, 229, 229, 229, 230, 230, 230, 229, 229, 229, 228, 229, 229, 229, 228, 231, 229, 228, 228, 230, 230, 230, 230, 230, 230, 230, 231, 231, 232, 231, 232, 233, 234, 234, 232, 232, 233, 235, 235, 235, 235, 236, 236, 236, 231, 212, 169, 121, 82, 70, 67, 65, 68, 74, 78, 81, 75, 76, 79, 77, 83, 80, 74, 70, 78, 96, 134, 159, 179, 193, 212, 221, 224, 222, 227, 226, 227, 226, 226, 228, 228, 228, 229, 228, 227, 228, 228, 228, 229, 228, 227, 227, 227, 226, 229, 227, 227, 228, 229, 227, 228, 228, 227, 227, 228, 229, 226, 226, 228, 229, 227, 228, 227, 226, 228, 228, 228, 226, 227, 223, 225, 228, 227, 224, 224, 227, 227, 227, 226, 225, 223, 222, 223, 225, 222, 218, 215, 213, 211, 208, 211, 212, 132, 209, 216, 211, 210, 214, 211, 209, 211, 212, 214, 213, 214, 216, 219, 219, 219, 218, 220, 219, 219, 219, 217, 219, 219, 219, 222, 221, 221, 222, 223, 222, 222, 222, 224, 222, 225, 224, 223, 225, 224, 227, 225, 225, 223, 225, 226, 226, 226, 225, 225, 228, 227, 226, 226, 226, 226, 227, 227, 227, 227, 227, 227, 228, 228, 226, 227, 226, 227, 226, 225, 226, 226, 227, 228, 227, 227, 227, 226, 228, 228, 226, 228, 227, 227, 229, 228, 227, 228, 228, 228, 229, 230, 227, 227, 228, 229, 228, 228, 228, 227, 230, 230, 230, 227, 229, 229, 230, 230, 228, 228, 227, 230, 230, 230, 229, 228, 230, 230, 229, 229, 228, 228, 230, 230, 229, 229, 229, 230, 231, 231, 229, 229, 229, 230, 231, 231, 230, 231, 231, 231, 234, 232, 232, 232, 233, 234, 234, 234, 234, 235, 236, 236, 237, 237, 236, 231, 215, 157, 89, 68, 69, 72, 78, 84, 86, 87, 88, 94, 94, 98, 111, 114, 123, 130, 118, 100, 88, 78, 69, 63, 63, 86, 115, 151, 175, 198, 214, 221, 226, 228, 226, 226, 227, 224, 228, 228, 229, 227, 227, 228, 228, 230, 228, 227, 227, 228, 228, 227, 228, 227, 228, 229, 229, 227, 228, 227, 227, 227, 228, 227, 224, 228, 229, 229, 229, 227, 228, 227, 227, 229, 227, 226, 225, 226, 226, 224, 227, 225, 227, 226, 227, 224, 223, 222, 223, 224, 226, 224, 218, 215, 205, 211, 210, 209, 212, 129, 208, 217, 212, 213, 212, 206, 207, 213, 215, 212, 215, 215, 219, 219, 218, 217, 218, 221, 219, 219, 218, 219, 218, 220, 221, 218, 221, 222, 221, 219, 223, 225, 222, 225, 226, 224, 224, 224, 224, 224, 228, 226, 226, 225, 224, 228, 226, 224, 224, 226, 229, 227, 228, 226, 226, 225, 228, 228, 228, 227, 227, 227, 228, 228, 226, 226, 227, 228, 227, 225, 225, 226, 226, 227, 227, 226, 228, 228, 228, 228, 227, 228, 227, 228, 227, 228, 227, 228, 228, 229, 229, 230, 228, 227, 228, 229, 228, 228, 228, 228, 229, 230, 229, 229, 229, 230, 230, 230, 229, 228, 227, 229, 229, 230, 229, 228, 228, 230, 230, 229, 229, 228, 231, 231, 229, 229, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 231, 232, 232, 232, 232, 232, 231, 232, 233, 233, 233, 233, 234, 234, 235, 236, 235, 232, 227, 203, 117, 73, 75, 96, 129, 147, 132, 103, 92, 102, 120, 146, 164, 181, 188, 200, 206, 210, 208, 207, 193, 168, 138, 93, 81, 73, 65, 72, 97, 127, 160, 198, 215, 226, 227, 227, 226, 226, 229, 229, 228, 227, 226, 227, 227, 230, 228, 227, 227, 227, 228, 229, 229, 229, 229, 228, 230, 229, 226, 226, 229, 229, 229, 226, 226, 227, 229, 228, 228, 229, 227, 227, 228, 226, 226, 224, 225, 227, 227, 226, 226, 222, 227, 225, 226, 225, 223, 224, 225, 226, 226, 224, 217, 213, 209, 210, 211, 209, 214, 124, 209, 216, 215, 215, 213, 215, 210, 216, 217, 217, 212, 217, 218, 220, 218, 218, 219, 219, 219, 219, 218, 222, 220, 219, 220, 216, 220, 221, 223, 222, 224, 224, 224, 226, 228, 226, 225, 224, 226, 227, 227, 227, 226, 224, 224, 226, 226, 224, 226, 226, 228, 226, 226, 226, 224, 224, 228, 229, 228, 227, 228, 227, 228, 227, 227, 225, 227, 229, 228, 226, 226, 225, 227, 224, 225, 225, 228, 227, 229, 228, 228, 227, 227, 228, 229, 228, 227, 226, 228, 229, 229, 229, 227, 228, 228, 229, 229, 229, 228, 228, 230, 230, 230, 230, 229, 230, 229, 228, 228, 228, 228, 230, 230, 230, 229, 229, 228, 229, 229, 229, 229, 229, 230, 231, 230, 229, 228, 230, 231, 231, 231, 230, 230, 231, 231, 231, 231, 230, 231, 232, 231, 231, 229, 230, 230, 232, 232, 233, 233, 232, 235, 234, 231, 224, 205, 110, 74, 86, 156, 201, 192, 146, 101, 105, 145, 178, 201, 215, 222, 226, 226, 224, 228, 229, 230, 230, 230, 228, 222, 209, 177, 125, 85, 77, 63, 78, 94, 116, 164, 206, 225, 226, 227, 226, 226, 229, 229, 228, 228, 228, 226, 227, 227, 227, 227, 228, 229, 229, 227, 228, 229, 229, 229, 229, 227, 227, 229, 229, 229, 228, 226, 228, 229, 229, 229, 228, 227, 227, 229, 227, 228, 224, 226, 227, 226, 228, 225, 224, 225, 224, 225, 224, 224, 224, 225, 226, 224, 223, 218, 213, 216, 211, 209, 210, 215, 141, 211, 216, 213, 217, 212, 212, 212, 215, 216, 218, 213, 217, 219, 217, 217, 219, 220, 219, 220, 222, 219, 220, 218, 219, 220, 217, 220, 222, 222, 223, 225, 224, 225, 227, 227, 226, 225, 222, 225, 227, 226, 226, 224, 224, 224, 225, 226, 226, 227, 226, 226, 229, 229, 227, 225, 226, 226, 228, 227, 227, 227, 227, 227, 228, 226, 227, 227, 228, 228, 227, 225, 226, 225, 228, 227, 226, 227, 227, 228, 229, 228, 228, 227, 228, 229, 229, 228, 227, 228, 229, 230, 230, 227, 228, 228, 229, 229, 229, 229, 229, 229, 230, 230, 229, 228, 230, 230, 230, 228, 228, 229, 230, 229, 230, 229, 228, 229, 230, 230, 228, 229, 229, 229, 230, 230, 229, 229, 229, 231, 231, 230, 230, 228, 230, 232, 231, 229, 230, 231, 232, 233, 230, 230, 230, 231, 232, 231, 232, 232, 233, 234, 232, 226, 213, 147, 82, 95, 182, 217, 204, 155, 104, 122, 176, 210, 223, 226, 230, 230, 230, 230, 228, 228, 228, 230, 229, 229, 232, 232, 231, 228, 217, 187, 125, 81, 71, 72, 89, 100, 139, 194, 218, 224, 226, 228, 229, 229, 228, 229, 225, 225, 225, 228, 228, 227, 228, 230, 230, 228, 228, 229, 230, 230, 229, 227, 228, 229, 229, 229, 227, 228, 227, 229, 229, 228, 229, 226, 227, 228, 228, 226, 226, 227, 227, 227, 225, 225, 225, 224, 223, 225, 226, 222, 225, 227, 225, 223, 223, 218, 212, 213, 213, 210, 210, 215, 128, 210, 215, 218, 218, 214, 208, 213, 215, 214, 212, 216, 215, 219, 218, 215, 218, 218, 224, 223, 223, 220, 218, 217, 222, 216, 219, 223, 224, 224, 225, 224, 223, 224, 224, 225, 227, 224, 224, 224, 226, 227, 226, 226, 224, 224, 226, 223, 225, 225, 225, 226, 229, 228, 228, 226, 226, 228, 228, 228, 228, 227, 228, 228, 228, 228, 226, 228, 228, 228, 228, 226, 226, 227, 227, 228, 226, 226, 227, 229, 229, 229, 227, 227, 227, 228, 228, 228, 228, 227, 229, 229, 229, 228, 228, 228, 229, 230, 229, 228, 228, 230, 230, 230, 229, 228, 230, 231, 230, 229, 229, 229, 230, 230, 230, 229, 229, 229, 229, 230, 229, 229, 228, 227, 228, 230, 229, 229, 230, 231, 232, 230, 229, 228, 231, 231, 231, 231, 230, 231, 232, 233, 232, 231, 231, 231, 231, 232, 232, 233, 233, 232, 228, 217, 191, 76, 83, 181, 220, 212, 167, 103, 119, 185, 222, 227, 229, 229, 231, 230, 231, 230, 229, 229, 228, 229, 229, 229, 232, 232, 234, 232, 232, 228, 213, 174, 97, 93, 76, 95, 97, 131, 186, 213, 226, 229, 229, 229, 229, 228, 228, 227, 226, 228, 228, 226, 228, 230, 229, 229, 228, 228, 230, 229, 228, 228, 228, 230, 229, 228, 228, 228, 228, 230, 229, 228, 228, 228, 229, 229, 229, 226, 224, 225, 228, 227, 225, 225, 224, 226, 226, 224, 225, 224, 220, 224, 226, 225, 222, 219, 213, 213, 213, 211, 212, 215, 140, 213, 214, 217, 218, 214, 212, 212, 214, 214, 213, 216, 214, 216, 218, 217, 216, 219, 222, 222, 220, 217, 217, 219, 218, 219, 220, 224, 223, 225, 223, 225, 224, 224, 226, 225, 227, 223, 226, 227, 228, 227, 227, 226, 225, 223, 227, 226, 224, 226, 226, 228, 229, 228, 228, 227, 226, 227, 229, 227, 228, 228, 227, 228, 229, 228, 227, 229, 229, 228, 227, 227, 227, 228, 227, 228, 227, 226, 227, 227, 228, 229, 227, 227, 228, 228, 230, 228, 227, 226, 229, 228, 229, 228, 228, 230, 230, 230, 229, 228, 228, 229, 230, 229, 230, 229, 230, 230, 230, 229, 229, 229, 230, 230, 230, 228, 228, 229, 229, 230, 227, 228, 229, 231, 230, 229, 229, 230, 231, 231, 231, 230, 230, 229, 231, 231, 231, 231, 230, 230, 233, 232, 231, 231, 230, 231, 232, 232, 233, 233, 233, 232, 225, 211, 141, 77, 130, 220, 217, 197, 121, 98, 168, 219, 228, 229, 227, 229, 229, 230, 228, 228, 229, 229, 228, 229, 230, 228, 230, 231, 232, 231, 232, 232, 229, 221, 181, 109, 107, 92, 122, 109, 126, 195, 222, 227, 229, 229, 228, 228, 228, 226, 228, 228, 226, 227, 228, 228, 230, 228, 228, 228, 229, 229, 230, 228, 227, 230, 230, 230, 229, 227, 228, 230, 230, 228, 228, 227, 229, 228, 228, 227, 226, 226, 229, 227, 225, 224, 225, 226, 227, 224, 224, 221, 224, 225, 224, 227, 225, 220, 213, 215, 218, 211, 212, 215, 126, 211, 216, 218, 215, 214, 215, 212, 214, 216, 213, 215, 215, 218, 217, 218, 216, 218, 221, 224, 221, 219, 217, 221, 219, 220, 220, 222, 222, 224, 224, 223, 224, 223, 224, 224, 226, 222, 225, 225, 225, 227, 227, 226, 225, 225, 228, 226, 226, 227, 229, 228, 229, 229, 227, 226, 228, 228, 228, 227, 228, 227, 228, 228, 228, 227, 228, 228, 230, 229, 230, 228, 228, 229, 228, 227, 227, 227, 228, 226, 229, 228, 227, 227, 228, 228, 229, 228, 229, 228, 228, 229, 229, 228, 228, 229, 230, 230, 229, 228, 228, 229, 230, 230, 229, 229, 229, 229, 230, 229, 229, 229, 230, 231, 230, 229, 229, 230, 231, 230, 229, 228, 230, 230, 231, 231, 229, 230, 230, 231, 231, 230, 230, 229, 231, 232, 231, 231, 231, 232, 233, 232, 232, 232, 231, 232, 232, 233, 233, 233, 233, 230, 222, 209, 93, 78, 193, 222, 213, 168, 97, 123, 203, 226, 226, 227, 227, 230, 230, 230, 228, 226, 229, 229, 230, 230, 228, 228, 229, 231, 231, 231, 231, 231, 233, 229, 219, 173, 135, 101, 143, 126, 96, 152, 212, 227, 228, 229, 229, 228, 229, 228, 229, 228, 227, 226, 229, 229, 230, 229, 229, 228, 231, 229, 230, 228, 228, 230, 230, 231, 228, 228, 230, 230, 229, 228, 228, 228, 229, 228, 227, 226, 225, 224, 227, 229, 228, 225, 226, 227, 225, 224, 225, 221, 221, 224, 225, 226, 224, 221, 213, 217, 219, 216, 215, 217, 121, 211, 217, 218, 214, 215, 216, 218, 214, 218, 216, 219, 217, 216, 219, 220, 219, 220, 224, 224, 224, 222, 221, 221, 220, 221, 219, 224, 221, 225, 223, 224, 222, 222, 224, 222, 225, 223, 224, 224, 226, 227, 227, 226, 227, 227, 227, 228, 227, 227, 228, 230, 229, 229, 227, 227, 229, 230, 228, 228, 227, 226, 227, 229, 228, 228, 227, 229, 229, 230, 230, 229, 228, 227, 228, 227, 226, 228, 227, 228, 226, 228, 227, 227, 228, 228, 228, 228, 228, 228, 229, 229, 229, 229, 229, 230, 230, 230, 228, 228, 229, 229, 229, 229, 229, 229, 229, 230, 230, 228, 229, 229, 230, 231, 230, 230, 229, 229, 231, 230, 228, 229, 229, 230, 231, 231, 230, 231, 231, 232, 232, 229, 228, 230, 230, 231, 230, 230, 231, 231, 233, 232, 232, 231, 231, 232, 233, 233, 231, 232, 232, 228, 219, 196, 94, 102, 216, 221, 211, 133, 94, 157, 218, 228, 227, 228, 228, 230, 230, 229, 226, 228, 227, 230, 229, 229, 228, 228, 229, 229, 228, 231, 232, 231, 232, 229, 227, 216, 137, 170, 114, 163, 107, 99, 189, 224, 229, 230, 228, 227, 229, 229, 229, 229, 227, 228, 229, 229, 229, 229, 229, 228, 231, 229, 229, 228, 228, 229, 230, 230, 227, 229, 229, 230, 229, 228, 229, 228, 228, 228, 227, 227, 226, 224, 226, 228, 228, 226, 227, 227, 226, 226, 224, 221, 222, 225, 225, 225, 223, 221, 218, 218, 216, 214, 214, 219, 132, 213, 219, 220, 217, 215, 217, 217, 213, 216, 216, 215, 220, 217, 220, 221, 219, 219, 224, 225, 220, 220, 221, 220, 220, 221, 219, 221, 222, 225, 223, 225, 223, 224, 225, 223, 224, 223, 225, 225, 227, 228, 226, 226, 224, 225, 226, 226, 226, 227, 228, 229, 229, 229, 228, 227, 227, 228, 229, 229, 227, 228, 227, 229, 230, 228, 227, 229, 230, 229, 227, 228, 228, 228, 229, 229, 227, 226, 228, 228, 228, 228, 227, 227, 229, 229, 229, 229, 229, 228, 230, 230, 230, 228, 228, 230, 230, 231, 230, 229, 228, 230, 229, 229, 229, 229, 229, 230, 231, 229, 229, 230, 231, 231, 230, 229, 230, 229, 229, 229, 229, 229, 229, 230, 231, 231, 230, 230, 231, 232, 232, 230, 229, 229, 230, 231, 231, 230, 231, 232, 233, 233, 232, 231, 232, 232, 232, 233, 232, 232, 231, 227, 219, 175, 119, 136, 223, 219, 199, 108, 92, 184, 224, 227, 228, 227, 227, 229, 230, 229, 228, 226, 226, 226, 229, 229, 228, 226, 229, 230, 228, 230, 228, 231, 231, 230, 230, 221, 203, 186, 159, 178, 142, 81, 140, 216, 228, 229, 228, 228, 228, 229, 230, 229, 227, 228, 230, 231, 230, 229, 229, 229, 230, 229, 226, 228, 229, 229, 230, 231, 228, 228, 228, 230, 229, 230, 229, 229, 229, 229, 226, 226, 227, 226, 228, 228, 229, 227, 227, 227, 224, 225, 224, 221, 220, 223, 225, 226, 224, 221, 217, 218, 216, 216, 213, 218, 124, 215, 220, 221, 217, 215, 214, 217, 215, 214, 215, 215, 219, 218, 219, 220, 220, 221, 223, 224, 222, 219, 218, 220, 221, 224, 222, 220, 222, 225, 224, 224, 222, 221, 224, 223, 225, 223, 226, 225, 228, 228, 227, 224, 226, 224, 228, 226, 228, 227, 228, 228, 230, 229, 228, 228, 228, 229, 229, 227, 226, 228, 229, 229, 230, 229, 228, 229, 230, 230, 229, 227, 228, 228, 229, 229, 228, 228, 228, 228, 228, 228, 227, 227, 227, 229, 229, 227, 228, 228, 230, 230, 229, 228, 228, 230, 229, 230, 229, 229, 228, 230, 230, 229, 229, 229, 229, 230, 229, 229, 229, 229, 231, 231, 230, 229, 229, 229, 230, 230, 230, 230, 229, 230, 231, 231, 230, 231, 230, 232, 231, 230, 229, 230, 231, 231, 232, 230, 231, 231, 233, 233, 232, 231, 232, 233, 232, 233, 232, 232, 230, 227, 219, 166, 116, 159, 224, 217, 190, 99, 102, 202, 226, 228, 228, 226, 225, 227, 229, 227, 227, 227, 225, 226, 229, 229, 228, 227, 229, 230, 230, 228, 230, 230, 231, 230, 230, 227, 224, 180, 220, 157, 174, 95, 101, 205, 228, 228, 229, 229, 227, 228, 230, 227, 228, 228, 229, 230, 230, 228, 228, 229, 230, 229, 228, 229, 228, 230, 230, 230, 228, 228, 229, 231, 230, 229, 228, 228, 230, 229, 228, 225, 225, 226, 227, 227, 227, 228, 227, 228, 228, 227, 224, 222, 224, 224, 227, 226, 224, 221, 215, 217, 218, 217, 213, 219, 119, 213, 219, 221, 218, 217, 213, 216, 217, 215, 216, 216, 218, 221, 220, 220, 222, 222, 224, 221, 223, 222, 218, 218, 220, 222, 223, 221, 223, 224, 224, 221, 223, 222, 224, 225, 226, 224, 224, 225, 228, 227, 228, 225, 226, 227, 227, 228, 226, 226, 228, 230, 229, 230, 229, 227, 228, 229, 228, 227, 227, 227, 229, 229, 230, 229, 228, 229, 230, 229, 229, 227, 228, 227, 230, 229, 229, 228, 228, 230, 229, 230, 228, 228, 228, 230, 230, 229, 229, 229, 229, 230, 229, 229, 228, 229, 229, 229, 229, 229, 228, 230, 230, 229, 229, 229, 228, 229, 230, 230, 229, 229, 230, 231, 230, 230, 229, 230, 231, 231, 230, 229, 229, 230, 230, 230, 230, 230, 231, 232, 231, 230, 229, 230, 231, 231, 231, 229, 231, 231, 233, 232, 231, 230, 232, 233, 233, 233, 231, 231, 230, 228, 219, 152, 119, 178, 223, 214, 175, 93, 122, 211, 228, 226, 227, 228, 227, 226, 229, 228, 227, 228, 225, 227, 230, 229, 229, 230, 229, 230, 229, 228, 230, 230, 230, 231, 228, 229, 226, 193, 226, 166, 193, 116, 79, 180, 226, 228, 225, 227, 228, 228, 229, 227, 229, 229, 230, 229, 230, 229, 228, 229, 230, 229, 229, 229, 229, 229, 229, 230, 229, 228, 230, 230, 230, 229, 227, 229, 230, 230, 229, 225, 224, 226, 228, 228, 227, 229, 228, 228, 227, 226, 225, 223, 226, 226, 227, 226, 226, 223, 216, 216, 217, 216, 212, 218, 118, 214, 218, 220, 215, 218, 216, 215, 221, 216, 215, 217, 219, 221, 221, 222, 224, 225, 220, 224, 222, 224, 218, 221, 224, 223, 223, 221, 224, 224, 224, 223, 223, 223, 224, 223, 225, 223, 223, 226, 226, 228, 228, 225, 227, 227, 227, 228, 226, 226, 228, 230, 230, 229, 228, 227, 229, 230, 228, 228, 228, 228, 229, 230, 230, 228, 228, 230, 229, 229, 229, 228, 228, 228, 229, 228, 228, 228, 228, 230, 230, 230, 228, 228, 229, 230, 228, 228, 229, 229, 229, 230, 230, 229, 228, 229, 229, 229, 229, 229, 229, 230, 230, 229, 229, 229, 230, 230, 230, 230, 230, 230, 230, 230, 230, 230, 229, 230, 230, 231, 228, 229, 229, 230, 230, 230, 229, 230, 231, 232, 231, 230, 229, 229, 231, 231, 232, 230, 231, 232, 232, 232, 231, 231, 231, 232, 233, 232, 232, 232, 230, 226, 223, 146, 129, 193, 224, 213, 163, 93, 135, 217, 228, 226, 226, 226, 226, 227, 228, 228, 227, 227, 226, 229, 230, 229, 230, 230, 230, 230, 229, 229, 229, 230, 230, 230, 229, 230, 223, 206, 214, 167, 197, 147, 78, 156, 223, 229, 226, 226, 227, 229, 229, 228, 228, 229, 230, 231, 230, 228, 228, 229, 231, 231, 230, 229, 230, 229, 230, 230, 229, 229, 229, 231, 230, 230, 230, 228, 230, 230, 229, 225, 226, 226, 228, 228, 228, 229, 227, 227, 228, 226, 225, 225, 225, 227, 225, 225, 227, 223, 215, 211, 218, 214, 214, 216, 135, 215, 217, 217, 216, 215, 215, 218, 215, 216, 216, 219, 223, 223, 223, 221, 221, 222, 221, 221, 222, 221, 223, 223, 224, 222, 223, 223, 222, 225, 224, 223, 221, 221, 224, 222, 223, 222, 224, 227, 227, 227, 228, 226, 226, 226, 228, 228, 228, 227, 228, 230, 230, 229, 228, 228, 227, 230, 230, 229, 228, 228, 230, 230, 230, 229, 229, 230, 230, 230, 229, 228, 228, 228, 227, 229, 229, 228, 228, 230, 229, 229, 229, 228, 229, 230, 229, 228, 228, 228, 229, 230, 230, 229, 229, 230, 230, 230, 229, 229, 229, 231, 230, 230, 229, 230, 229, 230, 230, 229, 229, 230, 230, 230, 230, 230, 229, 230, 230, 231, 229, 229, 229, 230, 229, 230, 230, 230, 230, 231, 232, 231, 230, 231, 231, 230, 231, 230, 231, 232, 232, 232, 231, 231, 231, 232, 232, 232, 230, 231, 230, 224, 222, 139, 126, 201, 221, 214, 152, 85, 148, 219, 228, 228, 227, 227, 225, 228, 227, 227, 229, 226, 226, 229, 229, 229, 230, 230, 229, 230, 230, 229, 229, 229, 230, 228, 230, 230, 221, 219, 179, 165, 189, 169, 75, 124, 214, 227, 225, 226, 226, 229, 226, 225, 229, 229, 230, 230, 230, 229, 228, 228, 230, 230, 230, 229, 230, 230, 231, 231, 229, 229, 229, 230, 230, 230, 229, 229, 230, 230, 228, 227, 226, 226, 228, 228, 230, 227, 228, 227, 229, 229, 227, 227, 227, 228, 226, 225, 227, 222, 216, 213, 218, 218, 212, 219, 133, 215, 216, 215, 214, 213, 213, 215, 220, 217, 216, 220, 223, 223, 224, 223, 221, 221, 223, 222, 222, 222, 222, 222, 219, 224, 221, 223, 223, 226, 222, 223, 222, 220, 224, 220, 222, 223, 224, 227, 228, 227, 229, 228, 228, 225, 227, 228, 228, 227, 228, 229, 231, 229, 228, 228, 228, 230, 229, 228, 229, 227, 230, 229, 229, 228, 229, 230, 230, 230, 229, 228, 228, 228, 230, 229, 228, 227, 229, 229, 230, 229, 228, 228, 229, 229, 229, 228, 229, 229, 230, 231, 230, 229, 228, 230, 229, 229, 229, 229, 229, 231, 231, 230, 229, 229, 229, 230, 230, 229, 228, 229, 230, 230, 230, 229, 229, 229, 231, 231, 229, 229, 230, 230, 230, 230, 230, 230, 230, 230, 230, 230, 230, 230, 231, 231, 231, 230, 230, 232, 232, 233, 232, 231, 231, 231, 232, 232, 231, 230, 229, 224, 221, 135, 119, 202, 222, 214, 145, 85, 152, 219, 228, 230, 226, 227, 227, 228, 227, 229, 229, 229, 227, 229, 230, 231, 229, 228, 229, 230, 230, 230, 229, 228, 227, 229, 229, 228, 223, 226, 169, 191, 180, 185, 84, 104, 212, 228, 225, 225, 227, 229, 225, 227, 228, 229, 231, 230, 230, 229, 227, 230, 230, 231, 230, 230, 230, 230, 229, 231, 228, 228, 229, 230, 229, 229, 227, 229, 229, 229, 229, 228, 229, 227, 229, 227, 229, 228, 229, 228, 230, 229, 228, 227, 226, 226, 228, 226, 228, 223, 214, 214, 218, 215, 212, 220, 136, 215, 218, 216, 215, 214, 216, 216, 220, 219, 218, 218, 223, 222, 224, 222, 221, 223, 222, 222, 223, 224, 222, 223, 220, 224, 225, 223, 223, 226, 224, 224, 224, 221, 224, 221, 222, 223, 224, 227, 226, 228, 229, 227, 227, 226, 228, 230, 229, 228, 229, 229, 230, 229, 229, 228, 228, 228, 229, 229, 228, 229, 230, 229, 229, 229, 229, 229, 230, 230, 229, 229, 228, 229, 230, 229, 228, 227, 229, 230, 229, 229, 228, 228, 229, 230, 230, 229, 229, 229, 230, 231, 230, 229, 229, 229, 230, 230, 229, 229, 229, 230, 230, 230, 230, 230, 230, 230, 230, 229, 229, 228, 231, 230, 230, 229, 230, 230, 230, 231, 229, 229, 229, 230, 231, 230, 229, 230, 230, 230, 231, 231, 230, 230, 232, 232, 231, 231, 231, 232, 232, 233, 232, 232, 230, 229, 223, 228, 231, 231, 228, 223, 212, 122, 108, 213, 219, 210, 142, 81, 166, 222, 228, 229, 226, 228, 227, 228, 228, 228, 228, 228, 225, 229, 230, 230, 230, 230, 230, 230, 231, 229, 229, 227, 228, 225, 229, 226, 227, 226, 166, 202, 168, 191, 97, 94, 205, 226, 225, 224, 224, 226, 228, 227, 227, 227, 229, 231, 231, 229, 228, 229, 230, 230, 229, 229, 229, 230, 230, 229, 229, 229, 228, 229, 228, 230, 229, 228, 229, 229, 230, 228, 228, 229, 229, 228, 229, 227, 228, 229, 230, 228, 227, 227, 226, 227, 226, 228, 225, 223, 217, 216, 219, 215, 211, 219, 126, 215, 218, 217, 216, 215, 216, 218, 220, 219, 216, 221, 224, 222, 225, 219, 220, 223, 223, 220, 222, 222, 224, 222, 223, 225, 224, 222, 224, 228, 226, 224, 222, 222, 224, 223, 225, 225, 227, 227, 227, 228, 229, 227, 228, 228, 229, 230, 228, 229, 229, 230, 230, 229, 229, 228, 230, 230, 230, 229, 228, 229, 230, 230, 231, 228, 228, 228, 230, 231, 230, 229, 229, 229, 230, 228, 228, 227, 228, 230, 230, 229, 229, 229, 229, 230, 230, 229, 229, 229, 231, 230, 230, 229, 229, 230, 230, 230, 229, 229, 230, 230, 231, 230, 229, 229, 230, 230, 230, 228, 229, 229, 231, 231, 230, 230, 229, 230, 231, 231, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 232, 230, 230, 231, 232, 233, 232, 232, 233, 233, 234, 234, 232, 228, 223, 182, 124, 184, 229, 230, 226, 214, 178, 107, 110, 218, 219, 204, 145, 135, 162, 188, 198, 209, 216, 221, 219, 221, 225, 225, 227, 228, 229, 230, 229, 230, 230, 229, 230, 231, 231, 229, 228, 228, 228, 229, 227, 226, 226, 225, 163, 189, 162, 195, 105, 80, 200, 225, 222, 225, 224, 227, 228, 227, 228, 228, 229, 230, 230, 230, 228, 230, 230, 230, 230, 230, 229, 229, 229, 230, 228, 229, 227, 229, 229, 230, 228, 228, 227, 228, 229, 228, 228, 229, 230, 229, 229, 228, 228, 229, 230, 229, 228, 227, 227, 229, 227, 226, 225, 223, 218, 216, 218, 219, 215, 221, 131, 215, 220, 215, 216, 217, 217, 217, 222, 220, 219, 220, 221, 223, 224, 219, 222, 221, 222, 222, 222, 221, 226, 223, 224, 224, 221, 224, 223, 228, 227, 227, 224, 224, 225, 223, 225, 224, 225, 227, 228, 228, 228, 228, 228, 227, 230, 230, 229, 228, 229, 230, 230, 231, 229, 229, 229, 229, 230, 229, 228, 229, 230, 230, 229, 228, 229, 230, 231, 230, 229, 227, 227, 229, 229, 229, 228, 228, 229, 230, 230, 229, 228, 229, 230, 230, 230, 229, 228, 229, 230, 231, 230, 229, 229, 230, 230, 230, 229, 229, 230, 231, 231, 230, 230, 229, 230, 231, 231, 229, 229, 229, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 232, 231, 231, 231, 231, 232, 232, 231, 231, 231, 233, 234, 233, 233, 234, 235, 235, 236, 232, 228, 221, 128, 129, 113, 223, 226, 213, 175, 119, 92, 151, 203, 185, 160, 148, 147, 136, 140, 136, 137, 146, 170, 179, 183, 193, 199, 210, 222, 227, 228, 229, 229, 230, 230, 229, 231, 231, 229, 226, 223, 219, 214, 213, 213, 217, 216, 173, 208, 146, 194, 110, 76, 183, 222, 225, 226, 227, 227, 228, 226, 228, 229, 230, 229, 229, 228, 228, 229, 230, 231, 230, 230, 230, 230, 230, 230, 229, 230, 223, 229, 230, 229, 228, 229, 228, 229, 229, 228, 227, 228, 229, 229, 229, 228, 228, 228, 230, 228, 228, 228, 227, 227, 227, 226, 227, 223, 221, 220, 216, 215, 214, 220, 133, 214, 219, 216, 221, 213, 219, 218, 219, 222, 221, 220, 221, 220, 223, 223, 222, 221, 221, 221, 221, 224, 225, 221, 223, 226, 223, 225, 225, 226, 226, 226, 224, 224, 225, 224, 226, 226, 225, 227, 229, 229, 227, 227, 227, 227, 230, 229, 229, 226, 229, 230, 230, 231, 229, 229, 230, 229, 230, 229, 228, 228, 230, 230, 230, 229, 229, 229, 230, 230, 229, 229, 228, 229, 229, 229, 229, 229, 228, 230, 230, 229, 228, 229, 230, 230, 230, 229, 229, 229, 230, 231, 230, 229, 230, 230, 230, 230, 229, 229, 230, 231, 231, 230, 230, 229, 230, 231, 231, 230, 230, 230, 230, 231, 230, 230, 229, 230, 232, 230, 231, 231, 231, 232, 232, 232, 232, 231, 231, 232, 232, 231, 232, 232, 233, 234, 234, 234, 234, 235, 237, 237, 235, 231, 222, 172, 111, 113, 193, 215, 197, 139, 100, 103, 132, 139, 130, 133, 130, 134, 120, 120, 124, 115, 115, 118, 132, 137, 116, 131, 154, 189, 212, 224, 231, 230, 232, 232, 233, 232, 230, 217, 191, 173, 155, 150, 143, 135, 140, 139, 126, 198, 121, 164, 91, 104, 168, 219, 223, 224, 227, 227, 227, 227, 228, 227, 229, 229, 229, 228, 227, 228, 230, 231, 229, 229, 230, 231, 231, 231, 230, 229, 227, 230, 231, 229, 229, 229, 229, 230, 230, 229, 228, 229, 230, 229, 230, 229, 228, 229, 229, 226, 228, 227, 228, 229, 226, 226, 225, 221, 220, 220, 217, 215, 212, 218, 124, 214, 219, 220, 216, 219, 219, 223, 218, 222, 220, 220, 221, 224, 224, 221, 223, 223, 224, 221, 221, 223, 224, 218, 224, 226, 223, 224, 225, 227, 227, 226, 224, 225, 224, 225, 226, 225, 226, 227, 228, 229, 228, 228, 228, 229, 230, 230, 227, 227, 229, 230, 230, 228, 230, 228, 229, 229, 230, 229, 229, 229, 230, 231, 230, 229, 229, 230, 231, 230, 229, 229, 228, 229, 230, 230, 228, 228, 229, 230, 230, 229, 229, 229, 230, 230, 229, 229, 230, 230, 230, 231, 230, 230, 229, 230, 230, 230, 229, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 229, 231, 231, 231, 231, 230, 231, 232, 232, 232, 231, 231, 231, 232, 233, 233, 232, 232, 234, 235, 234, 234, 234, 235, 237, 237, 237, 235, 231, 222, 148, 135, 107, 137, 127, 99, 125, 134, 131, 127, 126, 124, 123, 128, 127, 124, 129, 130, 123, 122, 116, 128, 120, 83, 87, 113, 163, 199, 227, 232, 232, 232, 231, 224, 197, 168, 155, 153, 141, 145, 139, 134, 137, 134, 129, 127, 117, 120, 111, 101, 114, 173, 158, 186, 220, 216, 214, 225, 229, 228, 229, 229, 229, 228, 227, 229, 229, 230, 229, 228, 230, 230, 230, 231, 229, 229, 230, 231, 231, 230, 230, 230, 230, 230, 230, 229, 229, 228, 230, 230, 228, 228, 228, 228, 229, 228, 227, 226, 227, 226, 226, 225, 224, 220, 219, 218, 220, 216, 216, 217, 122, 210, 217, 221, 220, 217, 217, 219, 216, 220, 222, 219, 224, 222, 224, 222, 221, 224, 222, 222, 224, 223, 224, 222, 221, 224, 223, 222, 225, 228, 227, 226, 226, 225, 226, 227, 228, 225, 225, 226, 228, 228, 229, 229, 229, 228, 231, 230, 227, 228, 230, 231, 231, 230, 230, 229, 228, 229, 231, 230, 229, 230, 230, 230, 230, 230, 229, 229, 230, 230, 229, 229, 229, 229, 229, 230, 228, 229, 229, 229, 229, 229, 229, 229, 230, 230, 229, 229, 229, 229, 230, 230, 230, 229, 229, 230, 230, 231, 230, 230, 229, 231, 231, 230, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 231, 231, 230, 232, 232, 232, 231, 231, 231, 232, 232, 232, 232, 232, 233, 234, 234, 234, 234, 234, 235, 237, 237, 234, 232, 227, 159, 156, 123, 99, 123, 133, 139, 145, 140, 138, 142, 136, 142, 136, 138, 140, 142, 134, 131, 122, 122, 124, 128, 103, 64, 67, 93, 147, 202, 229, 231, 228, 221, 185, 162, 162, 156, 162, 161, 160, 162, 152, 155, 147, 149, 137, 127, 117, 114, 125, 128, 107, 128, 86, 163, 132, 131, 199, 226, 228, 228, 229, 229, 228, 227, 230, 230, 230, 229, 230, 230, 230, 231, 230, 229, 230, 229, 230, 231, 231, 230, 229, 230, 231, 230, 228, 228, 228, 230, 230, 228, 227, 228, 226, 228, 226, 227, 225, 223, 226, 225, 223, 223, 220, 217, 218, 220, 219, 212, 218, 116, 211, 217, 218, 218, 217, 217, 216, 218, 217, 220, 218, 221, 224, 223, 222, 220, 223, 220, 224, 226, 224, 223, 222, 221, 223, 222, 223, 223, 226, 227, 226, 225, 226, 224, 227, 225, 226, 227, 227, 227, 228, 229, 228, 229, 230, 231, 230, 228, 229, 230, 230, 231, 230, 230, 229, 230, 229, 230, 229, 229, 228, 230, 230, 230, 229, 229, 230, 230, 230, 230, 229, 228, 228, 229, 227, 229, 229, 229, 229, 229, 229, 228, 229, 230, 230, 230, 229, 229, 228, 229, 230, 230, 229, 229, 230, 230, 230, 230, 230, 229, 230, 231, 231, 229, 230, 230, 231, 231, 230, 230, 229, 231, 231, 231, 230, 231, 231, 232, 232, 231, 231, 231, 231, 233, 231, 230, 231, 231, 232, 233, 233, 232, 232, 233, 234, 234, 234, 234, 235, 235, 236, 236, 234, 230, 222, 163, 130, 111, 133, 135, 141, 148, 145, 139, 137, 144, 143, 148, 148, 145, 148, 147, 146, 141, 133, 131, 127, 124, 130, 77, 70, 92, 104, 160, 212, 223, 219, 180, 151, 136, 135, 127, 137, 158, 160, 163, 168, 168, 164, 165, 157, 152, 142, 131, 132, 126, 128, 116, 84, 70, 64, 78, 174, 225, 227, 229, 228, 230, 227, 227, 228, 229, 230, 230, 230, 230, 231, 230, 230, 230, 229, 229, 231, 230, 231, 229, 230, 231, 230, 229, 229, 229, 229, 230, 229, 229, 227, 226, 226, 228, 229, 227, 227, 225, 228, 227, 223, 224, 218, 218, 219, 216, 218, 216, 219, 135, 213, 221, 220, 220, 218, 220, 217, 220, 218, 215, 219, 219, 224, 224, 221, 222, 223, 224, 224, 227, 226, 224, 224, 224, 226, 224, 224, 224, 227, 227, 226, 226, 225, 224, 225, 227, 226, 226, 227, 229, 229, 230, 228, 228, 229, 231, 230, 230, 228, 229, 229, 230, 231, 229, 229, 229, 230, 230, 230, 229, 228, 230, 230, 230, 229, 229, 230, 231, 230, 230, 228, 229, 229, 227, 229, 229, 228, 229, 230, 230, 230, 229, 228, 230, 230, 230, 229, 229, 228, 230, 230, 230, 229, 229, 230, 231, 231, 230, 230, 229, 231, 231, 231, 230, 229, 230, 232, 232, 231, 230, 230, 231, 231, 231, 230, 230, 231, 231, 232, 231, 231, 231, 232, 231, 232, 231, 232, 232, 233, 234, 233, 232, 232, 233, 235, 235, 235, 234, 235, 236, 237, 236, 233, 228, 213, 143, 141, 120, 119, 129, 145, 145, 147, 148, 150, 153, 153, 164, 161, 162, 160, 163, 155, 150, 144, 137, 125, 134, 129, 96, 66, 109, 86, 113, 140, 163, 157, 102, 60, 54, 54, 58, 71, 90, 106, 143, 162, 167, 174, 173, 169, 165, 158, 148, 144, 137, 128, 112, 104, 84, 57, 79, 153, 206, 221, 227, 229, 230, 228, 227, 228, 229, 230, 231, 230, 229, 230, 230, 231, 230, 229, 229, 230, 230, 231, 229, 230, 230, 229, 229, 229, 229, 229, 230, 229, 230, 229, 228, 226, 228, 226, 228, 227, 226, 226, 226, 226, 224, 219, 219, 218, 220, 219, 218, 221, 148, 215, 220, 219, 219, 219, 219, 220, 220, 221, 217, 217, 220, 222, 222, 224, 222, 223, 224, 226, 226, 227, 224, 222, 225, 226, 224, 225, 226, 224, 226, 227, 227, 225, 225, 227, 225, 228, 227, 226, 227, 229, 229, 228, 227, 228, 230, 231, 230, 228, 228, 230, 230, 230, 230, 230, 229, 231, 231, 230, 229, 230, 231, 231, 230, 229, 229, 230, 230, 231, 230, 229, 229, 229, 230, 228, 229, 228, 228, 230, 231, 230, 229, 229, 229, 231, 231, 229, 228, 229, 230, 230, 231, 229, 229, 229, 230, 230, 230, 229, 229, 231, 231, 231, 230, 229, 230, 231, 232, 231, 230, 230, 231, 231, 231, 231, 230, 231, 231, 232, 231, 230, 230, 232, 231, 231, 231, 231, 231, 232, 233, 232, 232, 232, 233, 234, 234, 234, 234, 235, 236, 236, 234, 229, 217, 190, 144, 135, 124, 130, 136, 144, 147, 154, 158, 163, 165, 169, 170, 168, 171, 169, 172, 166, 167, 158, 143, 133, 129, 86, 103, 55, 126, 92, 148, 107, 100, 85, 42, 51, 57, 63, 64, 60, 53, 53, 63, 77, 110, 155, 175, 170, 172, 177, 170, 165, 154, 150, 132, 123, 110, 111, 75, 85, 143, 188, 217, 228, 228, 227, 227, 228, 229, 231, 230, 230, 230, 230, 230, 230, 230, 229, 228, 229, 229, 230, 230, 229, 230, 230, 229, 229, 230, 229, 229, 230, 229, 227, 227, 227, 227, 227, 227, 227, 226, 228, 229, 228, 225, 224, 219, 215, 220, 219, 217, 223, 130, 215, 222, 220, 220, 221, 220, 221, 222, 221, 220, 221, 222, 224, 226, 225, 222, 223, 224, 224, 224, 225, 224, 222, 225, 225, 225, 225, 225, 225, 226, 226, 227, 226, 226, 228, 227, 227, 228, 226, 227, 229, 229, 227, 226, 228, 230, 231, 229, 229, 228, 230, 230, 230, 229, 230, 230, 231, 231, 230, 229, 230, 231, 231, 230, 229, 229, 229, 231, 231, 229, 229, 229, 230, 229, 230, 228, 228, 228, 230, 231, 230, 228, 228, 230, 230, 230, 230, 229, 229, 230, 231, 229, 229, 229, 230, 231, 231, 229, 229, 229, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 232, 231, 230, 230, 231, 232, 232, 231, 231, 232, 233, 233, 232, 232, 233, 234, 234, 234, 234, 234, 235, 236, 234, 228, 206, 174, 166, 153, 151, 143, 142, 151, 155, 152, 163, 168, 174, 173, 179, 178, 179, 176, 181, 174, 176, 172, 164, 149, 128, 90, 63, 72, 66, 67, 76, 140, 88, 159, 123, 43, 54, 76, 86, 77, 59, 58, 66, 57, 56, 78, 152, 113, 154, 174, 181, 186, 181, 173, 166, 158, 142, 123, 117, 115, 82, 66, 112, 173, 214, 223, 226, 227, 228, 229, 230, 230, 230, 230, 230, 231, 229, 229, 230, 229, 230, 230, 230, 230, 229, 229, 230, 229, 230, 230, 230, 230, 229, 229, 228, 228, 228, 229, 227, 228, 226, 227, 227, 226, 228, 228, 225, 220, 216, 221, 221, 215, 219, 137, 218, 223, 224, 221, 221, 219, 224, 221, 219, 222, 220, 223, 226, 227, 225, 225, 226, 226, 224, 223, 223, 224, 224, 227, 225, 225, 225, 224, 227, 225, 226, 227, 224, 227, 227, 228, 228, 227, 226, 228, 230, 228, 228, 227, 229, 229, 230, 229, 230, 229, 229, 230, 230, 229, 230, 230, 230, 230, 230, 229, 229, 231, 230, 230, 229, 229, 230, 231, 230, 229, 228, 229, 228, 230, 230, 229, 228, 229, 230, 230, 230, 229, 229, 230, 231, 230, 229, 229, 229, 230, 230, 230, 229, 229, 230, 231, 230, 229, 229, 230, 230, 231, 231, 230, 229, 231, 232, 231, 230, 230, 230, 232, 231, 231, 231, 230, 231, 232, 232, 231, 231, 230, 232, 232, 232, 231, 231, 232, 232, 233, 233, 232, 233, 234, 234, 235, 234, 235, 234, 233, 225, 195, 171, 157, 152, 144, 146, 146, 152, 158, 164, 169, 176, 173, 179, 184, 187, 187, 182, 182, 183, 190, 184, 180, 161, 136, 79, 54, 55, 59, 54, 64, 66, 108, 127, 87, 55, 44, 51, 76, 107, 136, 156, 149, 168, 160, 113, 162, 85, 57, 64, 112, 157, 185, 184, 181, 175, 171, 155, 148, 132, 112, 121, 75, 57, 97, 156, 208, 225, 227, 228, 230, 231, 231, 230, 230, 230, 230, 230, 225, 229, 230, 228, 231, 231, 230, 229, 229, 229, 230, 229, 229, 230, 230, 230, 230, 228, 229, 229, 229, 228, 226, 228, 227, 228, 227, 229, 226, 224, 222, 218, 222, 219, 219, 219, 150, 218, 222, 226, 220, 221, 220, 226, 223, 221, 223, 221, 223, 225, 223, 225, 226, 226, 225, 224, 225, 224, 224, 224, 224, 226, 224, 225, 226, 226, 226, 227, 225, 225, 227, 228, 229, 227, 226, 228, 230, 228, 229, 227, 226, 228, 229, 229, 228, 229, 229, 230, 231, 230, 230, 230, 230, 231, 230, 230, 230, 229, 229, 230, 230, 230, 229, 230, 231, 230, 230, 229, 229, 229, 230, 229, 228, 229, 229, 231, 230, 230, 229, 229, 230, 230, 230, 229, 230, 230, 231, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 232, 230, 230, 230, 231, 231, 232, 231, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 232, 233, 232, 233, 233, 233, 234, 235, 235, 234, 234, 230, 224, 188, 169, 156, 150, 151, 148, 155, 154, 163, 170, 178, 184, 183, 185, 187, 190, 192, 192, 188, 187, 188, 188, 184, 171, 135, 74, 57, 55, 57, 54, 63, 87, 109, 182, 210, 190, 65, 62, 71, 172, 185, 126, 144, 134, 160, 157, 139, 123, 50, 52, 53, 55, 71, 128, 171, 176, 180, 176, 166, 157, 143, 128, 123, 130, 70, 63, 93, 155, 208, 224, 229, 230, 231, 231, 230, 230, 230, 230, 229, 228, 225, 229, 226, 230, 230, 229, 229, 230, 229, 230, 229, 229, 230, 230, 230, 230, 226, 229, 229, 228, 229, 225, 228, 228, 229, 228, 228, 227, 225, 223, 221, 218, 219, 215, 222, 135, 219, 221, 224, 220, 221, 221, 222, 222, 220, 221, 221, 224, 225, 225, 225, 225, 226, 225, 224, 225, 225, 226, 225, 227, 226, 223, 225, 226, 226, 226, 227, 226, 224, 227, 229, 229, 228, 228, 228, 229, 227, 229, 228, 227, 227, 230, 230, 228, 228, 230, 231, 231, 230, 229, 229, 230, 231, 230, 229, 229, 229, 230, 230, 230, 230, 229, 230, 231, 231, 230, 229, 228, 230, 231, 228, 227, 229, 230, 231, 231, 230, 230, 230, 231, 230, 230, 229, 230, 229, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 231, 232, 231, 230, 230, 231, 232, 231, 231, 230, 231, 231, 231, 231, 230, 231, 231, 231, 231, 231, 231, 231, 232, 233, 232, 231, 231, 233, 233, 232, 233, 233, 233, 235, 234, 235, 233, 231, 223, 190, 168, 157, 150, 152, 152, 154, 162, 165, 174, 180, 188, 187, 193, 195, 195, 196, 192, 199, 196, 196, 192, 184, 171, 125, 64, 58, 58, 55, 57, 69, 97, 139, 139, 165, 182, 186, 114, 112, 146, 200, 106, 80, 60, 59, 65, 63, 61, 72, 67, 75, 66, 49, 61, 71, 86, 132, 166, 177, 179, 166, 161, 151, 130, 119, 117, 60, 70, 88, 156, 210, 226, 227, 230, 230, 229, 229, 230, 231, 230, 230, 224, 223, 230, 230, 230, 229, 229, 230, 230, 231, 229, 230, 229, 229, 229, 231, 229, 228, 230, 229, 228, 228, 229, 228, 228, 228, 228, 228, 226, 221, 219, 222, 220, 217, 222, 127, 216, 222, 223, 222, 222, 223, 222, 222, 219, 222, 219, 223, 225, 225, 224, 224, 225, 227, 225, 225, 224, 225, 224, 224, 226, 226, 227, 226, 226, 227, 227, 225, 225, 228, 228, 229, 228, 228, 229, 230, 230, 229, 228, 228, 229, 229, 230, 229, 229, 229, 231, 231, 230, 230, 229, 230, 231, 231, 229, 228, 229, 230, 230, 231, 230, 229, 230, 230, 230, 230, 228, 228, 230, 230, 229, 229, 229, 229, 230, 230, 230, 229, 229, 231, 230, 231, 229, 229, 230, 231, 231, 230, 230, 230, 230, 230, 231, 229, 229, 230, 231, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 231, 231, 230, 231, 231, 231, 231, 231, 232, 233, 232, 232, 232, 232, 232, 233, 233, 232, 233, 232, 235, 234, 234, 230, 225, 193, 168, 163, 156, 150, 152, 157, 165, 166, 174, 179, 185, 192, 195, 204, 200, 202, 201, 197, 201, 196, 191, 182, 156, 101, 68, 105, 153, 128, 99, 95, 107, 135, 134, 136, 143, 135, 142, 137, 136, 140, 139, 133, 125, 114, 105, 89, 71, 67, 69, 69, 79, 73, 67, 61, 55, 59, 56, 85, 151, 176, 173, 171, 163, 142, 123, 127, 110, 56, 60, 97, 175, 220, 228, 230, 229, 229, 229, 230, 232, 229, 229, 229, 230, 231, 230, 230, 229, 230, 231, 231, 231, 230, 229, 229, 231, 230, 230, 229, 228, 230, 231, 228, 228, 228, 225, 228, 230, 228, 227, 225, 221, 219, 222, 217, 217, 222, 126, 216, 222, 221, 220, 221, 221, 221, 221, 220, 220, 220, 222, 224, 225, 225, 222, 225, 226, 226, 227, 225, 226, 226, 224, 226, 226, 226, 226, 227, 228, 228, 225, 227, 228, 229, 230, 228, 227, 228, 229, 230, 230, 228, 227, 228, 229, 230, 229, 229, 230, 230, 230, 230, 229, 229, 230, 230, 230, 230, 228, 229, 230, 230, 231, 230, 230, 230, 231, 230, 229, 229, 229, 231, 231, 230, 229, 229, 229, 230, 230, 230, 230, 230, 230, 230, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 229, 229, 230, 231, 232, 231, 230, 229, 230, 231, 232, 230, 230, 230, 231, 231, 232, 230, 231, 231, 232, 232, 232, 231, 230, 232, 233, 233, 232, 231, 232, 233, 234, 232, 232, 234, 235, 234, 233, 228, 204, 169, 165, 160, 162, 159, 159, 164, 172, 176, 180, 185, 188, 200, 203, 208, 202, 207, 201, 203, 204, 193, 180, 145, 73, 60, 62, 86, 107, 100, 117, 131, 140, 145, 143, 147, 147, 149, 144, 141, 147, 147, 148, 145, 144, 151, 143, 132, 121, 108, 91, 81, 81, 76, 68, 66, 55, 51, 37, 51, 70, 137, 166, 176, 164, 148, 134, 121, 133, 83, 48, 75, 118, 195, 224, 229, 230, 230, 230, 230, 231, 231, 229, 229, 229, 231, 231, 230, 230, 229, 230, 231, 231, 230, 229, 229, 230, 230, 230, 229, 229, 230, 230, 230, 228, 228, 225, 228, 228, 227, 229, 225, 222, 220, 222, 218, 218, 222, 124, 217, 223, 223, 223, 219, 220, 220, 220, 217, 222, 221, 223, 226, 225, 224, 225, 225, 226, 228, 226, 224, 225, 225, 225, 225, 225, 225, 226, 227, 229, 227, 226, 227, 226, 229, 228, 228, 228, 228, 230, 230, 229, 229, 229, 229, 230, 231, 230, 230, 229, 230, 230, 230, 230, 229, 230, 231, 230, 229, 228, 229, 231, 231, 230, 230, 230, 230, 230, 230, 230, 230, 229, 230, 231, 231, 229, 229, 230, 231, 231, 231, 229, 230, 231, 231, 230, 229, 229, 230, 231, 231, 230, 229, 230, 231, 231, 230, 229, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 232, 232, 231, 230, 231, 231, 232, 232, 231, 232, 231, 232, 233, 233, 232, 232, 232, 233, 233, 233, 233, 233, 234, 234, 231, 220, 181, 163, 158, 163, 160, 166, 165, 174, 179, 183, 191, 195, 200, 210, 208, 221, 215, 214, 205, 203, 195, 169, 106, 64, 62, 66, 88, 106, 115, 133, 148, 153, 149, 145, 144, 150, 152, 156, 162, 165, 164, 168, 167, 176, 174, 179, 180, 173, 169, 159, 146, 123, 106, 87, 60, 61, 50, 48, 43, 49, 54, 68, 117, 162, 165, 161, 148, 126, 124, 130, 55, 52, 84, 146, 211, 228, 230, 228, 229, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 229, 229, 229, 230, 230, 229, 229, 230, 230, 231, 231, 230, 228, 228, 226, 226, 229, 227, 229, 225, 222, 219, 218, 218, 217, 224, 132, 216, 221, 225, 221, 221, 218, 219, 221, 220, 222, 221, 222, 225, 226, 224, 223, 225, 225, 225, 224, 222, 223, 224, 225, 224, 225, 225, 225, 228, 227, 228, 227, 226, 226, 229, 229, 228, 227, 229, 230, 230, 230, 230, 229, 229, 229, 230, 229, 229, 230, 230, 230, 230, 229, 230, 230, 231, 230, 230, 229, 230, 231, 230, 230, 230, 230, 229, 229, 230, 230, 229, 229, 230, 231, 231, 229, 229, 230, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 230, 230, 230, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 232, 231, 231, 231, 232, 233, 233, 232, 231, 232, 233, 233, 233, 233, 232, 234, 233, 229, 195, 172, 167, 164, 167, 166, 171, 176, 181, 189, 193, 193, 202, 206, 212, 233, 234, 220, 210, 204, 184, 143, 81, 67, 70, 83, 109, 120, 128, 147, 153, 150, 148, 145, 145, 155, 163, 162, 163, 171, 186, 191, 198, 200, 208, 210, 214, 218, 219, 210, 204, 192, 178, 168, 142, 111, 71, 51, 47, 51, 55, 54, 57, 68, 91, 152, 161, 156, 136, 123, 133, 83, 51, 65, 102, 192, 227, 229, 228, 229, 229, 231, 230, 230, 229, 229, 231, 231, 230, 230, 230, 230, 231, 230, 229, 228, 228, 231, 230, 230, 229, 230, 231, 231, 231, 229, 227, 226, 225, 228, 227, 229, 225, 224, 219, 220, 218, 218, 221, 138, 219, 224, 224, 221, 223, 220, 220, 220, 221, 222, 221, 225, 223, 224, 224, 224, 224, 225, 226, 223, 224, 224, 224, 225, 225, 226, 224, 226, 227, 226, 228, 227, 226, 227, 228, 228, 227, 228, 228, 229, 229, 229, 230, 228, 229, 230, 230, 229, 229, 230, 230, 230, 230, 229, 230, 229, 230, 230, 229, 229, 229, 230, 231, 230, 229, 229, 230, 230, 230, 230, 229, 229, 230, 230, 230, 229, 230, 230, 231, 230, 229, 229, 229, 230, 231, 231, 230, 230, 230, 230, 230, 230, 229, 230, 230, 231, 231, 229, 229, 229, 230, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 232, 232, 232, 231, 231, 230, 232, 232, 231, 231, 231, 233, 233, 233, 231, 231, 231, 234, 233, 233, 233, 233, 234, 231, 223, 182, 167, 164, 168, 168, 169, 176, 183, 188, 191, 197, 198, 205, 212, 224, 236, 234, 213, 198, 166, 105, 61, 60, 75, 108, 122, 133, 142, 150, 156, 148, 140, 147, 155, 160, 161, 166, 180, 189, 195, 200, 201, 204, 207, 206, 210, 217, 220, 226, 227, 229, 229, 225, 214, 195, 173, 150, 111, 67, 53, 57, 59, 61, 68, 65, 87, 145, 150, 149, 131, 124, 124, 48, 60, 74, 165, 220, 229, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 229, 230, 231, 231, 229, 227, 228, 229, 230, 230, 229, 230, 230, 230, 230, 229, 227, 226, 224, 226, 230, 228, 225, 223, 219, 220, 218, 216, 219, 124, 217, 224, 221, 223, 222, 222, 223, 224, 221, 222, 220, 223, 226, 224, 225, 226, 224, 225, 228, 225, 224, 224, 225, 225, 224, 224, 225, 225, 229, 226, 228, 227, 226, 228, 228, 228, 228, 228, 227, 229, 229, 230, 229, 228, 229, 230, 231, 229, 229, 229, 230, 231, 231, 230, 229, 228, 230, 229, 229, 228, 230, 231, 230, 230, 229, 230, 230, 230, 230, 230, 229, 229, 230, 231, 231, 229, 230, 229, 230, 230, 231, 230, 230, 230, 231, 231, 229, 230, 230, 231, 231, 230, 229, 229, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 230, 230, 230, 231, 232, 232, 231, 231, 231, 232, 233, 231, 231, 231, 233, 233, 232, 231, 231, 232, 233, 233, 233, 233, 232, 233, 229, 213, 175, 166, 167, 170, 173, 177, 181, 189, 186, 193, 199, 202, 210, 216, 221, 232, 220, 189, 125, 60, 53, 66, 99, 117, 126, 137, 152, 159, 154, 142, 142, 159, 160, 152, 156, 169, 178, 185, 194, 200, 196, 199, 202, 205, 207, 209, 213, 220, 224, 223, 226, 226, 229, 233, 232, 223, 205, 171, 145, 104, 54, 50, 62, 64, 68, 70, 84, 145, 144, 141, 121, 143, 55, 52, 81, 133, 214, 229, 228, 230, 231, 231, 232, 230, 230, 230, 231, 229, 231, 230, 229, 230, 230, 231, 230, 227, 227, 229, 230, 231, 229, 230, 230, 231, 229, 230, 228, 229, 226, 227, 230, 227, 222, 222, 218, 221, 222, 218, 217, 143, 217, 223, 224, 224, 222, 222, 223, 222, 223, 221, 221, 223, 225, 226, 225, 225, 226, 224, 227, 226, 222, 224, 224, 225, 224, 222, 224, 224, 226, 226, 229, 227, 227, 227, 229, 229, 229, 228, 228, 229, 230, 230, 228, 228, 230, 230, 230, 229, 229, 230, 231, 231, 231, 229, 229, 229, 229, 229, 229, 229, 230, 231, 230, 231, 229, 230, 230, 230, 230, 230, 229, 229, 230, 231, 230, 229, 229, 230, 230, 230, 230, 230, 230, 230, 231, 231, 229, 230, 230, 231, 231, 230, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 232, 230, 230, 230, 231, 232, 232, 231, 230, 232, 232, 232, 231, 231, 231, 232, 232, 233, 231, 232, 232, 234, 234, 234, 233, 233, 232, 229, 203, 174, 171, 172, 176, 177, 178, 186, 187, 193, 195, 203, 211, 209, 217, 213, 208, 166, 79, 64, 67, 88, 104, 121, 126, 147, 158, 156, 150, 142, 150, 165, 156, 152, 155, 174, 177, 178, 169, 161, 151, 141, 140, 143, 148, 157, 171, 187, 206, 219, 223, 223, 226, 228, 228, 233, 232, 233, 224, 201, 168, 132, 77, 56, 55, 61, 68, 71, 99, 141, 142, 135, 137, 70, 52, 70, 108, 204, 228, 229, 228, 230, 232, 231, 230, 230, 230, 231, 231, 230, 229, 229, 230, 231, 230, 230, 228, 228, 229, 230, 229, 229, 230, 230, 231, 229, 228, 228, 228, 226, 227, 227, 226, 224, 223, 218, 221, 221, 216, 219, 123, 214, 225, 224, 223, 220, 220, 226, 226, 222, 220, 222, 224, 225, 226, 226, 225, 224, 227, 227, 225, 224, 223, 227, 225, 225, 223, 224, 223, 227, 227, 227, 226, 228, 228, 228, 229, 228, 228, 228, 229, 230, 230, 229, 229, 230, 230, 229, 228, 228, 229, 230, 230, 231, 229, 228, 229, 230, 229, 229, 229, 229, 230, 231, 231, 230, 230, 230, 230, 230, 230, 230, 229, 230, 231, 230, 229, 229, 230, 231, 230, 230, 230, 230, 230, 231, 231, 229, 230, 230, 231, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 231, 232, 232, 232, 231, 231, 232, 232, 232, 232, 232, 231, 232, 233, 233, 231, 232, 233, 233, 234, 234, 233, 233, 233, 230, 202, 180, 178, 180, 179, 185, 184, 193, 193, 201, 205, 207, 212, 208, 197, 170, 118, 66, 69, 104, 95, 106, 122, 129, 148, 160, 167, 158, 138, 159, 165, 155, 152, 163, 154, 144, 134, 93, 65, 54, 48, 53, 59, 106, 149, 52, 53, 68, 95, 136, 173, 201, 219, 225, 230, 228, 231, 233, 235, 234, 222, 194, 154, 106, 55, 45, 57, 62, 62, 102, 136, 144, 142, 91, 49, 65, 90, 193, 226, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 230, 230, 230, 230, 229, 229, 230, 229, 230, 229, 230, 229, 230, 230, 229, 228, 228, 228, 227, 227, 227, 225, 223, 221, 222, 216, 218, 218, 110, 212, 224, 225, 223, 222, 222, 226, 225, 224, 225, 224, 225, 226, 223, 226, 224, 224, 229, 226, 226, 223, 224, 226, 227, 228, 226, 227, 225, 226, 228, 228, 226, 227, 228, 228, 229, 228, 227, 227, 230, 230, 230, 229, 229, 229, 231, 230, 229, 229, 229, 230, 231, 230, 230, 229, 230, 231, 230, 229, 229, 229, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 230, 230, 229, 230, 229, 231, 230, 230, 229, 230, 231, 231, 231, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 231, 232, 232, 232, 231, 231, 232, 233, 233, 232, 231, 231, 232, 233, 233, 232, 232, 233, 233, 234, 234, 234, 233, 233, 231, 207, 183, 180, 182, 187, 190, 196, 197, 198, 201, 207, 208, 196, 169, 118, 67, 70, 93, 83, 107, 133, 124, 135, 153, 165, 169, 160, 145, 164, 165, 143, 148, 152, 129, 116, 78, 44, 46, 48, 55, 96, 93, 75, 89, 117, 67, 64, 68, 47, 52, 60, 81, 140, 189, 215, 227, 229, 230, 235, 237, 235, 230, 210, 170, 121, 59, 46, 50, 57, 70, 122, 146, 145, 95, 53, 68, 92, 189, 226, 228, 229, 231, 231, 231, 230, 230, 230, 232, 231, 231, 230, 230, 230, 231, 230, 229, 229, 229, 230, 231, 231, 229, 230, 229, 230, 230, 229, 228, 228, 230, 228, 227, 230, 224, 224, 222, 220, 220, 218, 221, 120, 216, 226, 222, 222, 221, 224, 226, 224, 224, 225, 225, 225, 225, 225, 225, 225, 225, 228, 227, 226, 225, 226, 226, 227, 227, 226, 227, 225, 227, 229, 227, 227, 228, 229, 230, 229, 228, 227, 228, 230, 230, 230, 228, 228, 230, 231, 230, 229, 229, 229, 230, 230, 230, 230, 228, 228, 230, 231, 230, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 230, 230, 229, 230, 231, 230, 230, 230, 230, 230, 231, 229, 230, 230, 231, 231, 231, 230, 229, 229, 231, 231, 230, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 232, 231, 230, 230, 230, 232, 232, 232, 231, 231, 232, 233, 233, 231, 231, 231, 232, 233, 233, 232, 232, 233, 234, 234, 234, 234, 234, 234, 231, 215, 180, 184, 187, 193, 196, 203, 198, 207, 200, 193, 171, 118, 75, 76, 100, 123, 123, 107, 127, 131, 138, 159, 172, 176, 157, 146, 169, 160, 145, 139, 120, 86, 59, 59, 115, 45, 40, 50, 80, 160, 163, 133, 61, 128, 121, 75, 93, 119, 78, 45, 44, 56, 76, 122, 190, 223, 230, 233, 235, 235, 236, 232, 220, 181, 134, 70, 53, 59, 70, 80, 141, 152, 84, 45, 58, 88, 194, 226, 230, 229, 231, 231, 231, 230, 229, 231, 231, 231, 231, 230, 229, 230, 231, 231, 229, 229, 230, 230, 231, 230, 228, 228, 230, 231, 230, 227, 227, 229, 230, 229, 229, 229, 224, 223, 220, 221, 224, 218, 222, 124, 213, 226, 223, 220, 218, 224, 226, 223, 225, 224, 224, 224, 227, 225, 224, 224, 225, 227, 226, 226, 225, 228, 228, 227, 227, 225, 227, 226, 228, 228, 227, 227, 227, 228, 230, 229, 227, 227, 228, 230, 229, 230, 229, 229, 230, 231, 231, 229, 229, 229, 231, 230, 230, 230, 227, 229, 231, 230, 230, 230, 230, 231, 230, 231, 230, 230, 230, 230, 231, 230, 230, 230, 230, 231, 230, 230, 229, 229, 230, 231, 231, 230, 230, 231, 231, 231, 230, 229, 229, 230, 230, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 230, 231, 232, 232, 231, 231, 232, 233, 232, 232, 231, 232, 232, 233, 233, 232, 232, 233, 234, 235, 234, 234, 235, 235, 232, 226, 191, 186, 191, 198, 205, 206, 198, 189, 162, 119, 81, 91, 117, 133, 140, 144, 138, 136, 138, 140, 159, 176, 176, 162, 145, 172, 166, 133, 127, 99, 90, 55, 47, 48, 91, 107, 43, 43, 86, 152, 169, 145, 116, 158, 62, 45, 51, 124, 151, 61, 46, 46, 45, 57, 79, 144, 206, 230, 232, 235, 236, 235, 233, 223, 187, 139, 78, 51, 55, 61, 118, 150, 62, 46, 58, 97, 200, 227, 228, 229, 231, 232, 231, 229, 230, 230, 231, 231, 231, 229, 230, 230, 231, 231, 229, 228, 230, 231, 230, 230, 228, 227, 230, 230, 230, 230, 229, 230, 230, 230, 230, 230, 226, 223, 219, 225, 222, 220, 222, 119, 214, 223, 224, 222, 218, 221, 227, 223, 225, 224, 224, 225, 225, 225, 223, 227, 225, 227, 225, 224, 224, 225, 227, 226, 227, 227, 226, 226, 229, 228, 229, 227, 227, 229, 229, 229, 227, 225, 227, 230, 230, 230, 229, 230, 230, 231, 231, 228, 229, 229, 230, 231, 229, 229, 228, 229, 231, 230, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 230, 230, 229, 229, 230, 231, 230, 230, 229, 230, 231, 230, 230, 229, 230, 231, 231, 230, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 232, 231, 230, 232, 232, 232, 231, 231, 231, 233, 233, 233, 232, 232, 233, 234, 235, 235, 234, 234, 236, 235, 230, 208, 190, 196, 197, 194, 186, 149, 106, 90, 105, 129, 137, 136, 140, 144, 141, 136, 137, 142, 162, 180, 182, 171, 142, 172, 167, 130, 110, 96, 77, 175, 68, 45, 46, 54, 120, 84, 48, 87, 141, 170, 150, 144, 160, 50, 42, 53, 86, 157, 127, 36, 38, 40, 43, 52, 80, 126, 180, 224, 232, 235, 235, 235, 234, 225, 190, 144, 76, 46, 63, 98, 145, 50, 47, 61, 126, 213, 228, 229, 229, 231, 231, 230, 229, 229, 228, 230, 230, 230, 229, 230, 230, 230, 231, 228, 229, 230, 230, 230, 229, 228, 227, 229, 230, 229, 230, 230, 229, 230, 230, 228, 230, 224, 222, 217, 225, 222, 219, 222, 111, 213, 224, 224, 221, 221, 221, 224, 221, 225, 226, 223, 225, 228, 225, 225, 227, 227, 226, 226, 225, 224, 226, 227, 226, 226, 227, 226, 224, 229, 227, 228, 228, 227, 228, 229, 230, 227, 226, 227, 229, 231, 230, 229, 229, 230, 231, 230, 229, 230, 229, 230, 230, 230, 230, 229, 229, 230, 231, 230, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 229, 230, 230, 230, 230, 229, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 231, 231, 230, 232, 232, 232, 231, 231, 231, 232, 232, 231, 231, 232, 233, 233, 233, 232, 232, 233, 234, 235, 235, 235, 235, 236, 236, 234, 224, 203, 202, 179, 148, 126, 114, 126, 146, 150, 154, 149, 141, 143, 142, 144, 141, 131, 154, 183, 186, 181, 146, 169, 174, 139, 92, 59, 62, 81, 121, 116, 98, 51, 95, 108, 147, 59, 69, 126, 167, 152, 151, 154, 45, 39, 46, 73, 150, 149, 39, 36, 39, 53, 64, 101, 164, 75, 152, 219, 233, 233, 235, 235, 234, 225, 188, 135, 68, 59, 87, 108, 46, 50, 74, 176, 225, 228, 230, 229, 230, 231, 231, 229, 229, 230, 231, 231, 230, 230, 229, 231, 230, 231, 229, 229, 229, 230, 230, 229, 227, 228, 230, 230, 231, 230, 230, 228, 230, 230, 230, 229, 224, 220, 218, 227, 219, 220, 220, 117, 213, 224, 223, 224, 225, 223, 225, 223, 223, 225, 226, 226, 228, 225, 226, 226, 225, 226, 227, 227, 225, 226, 226, 227, 227, 227, 226, 225, 228, 228, 228, 228, 226, 227, 228, 227, 227, 227, 228, 230, 230, 230, 228, 228, 229, 230, 231, 230, 229, 230, 230, 230, 230, 229, 230, 230, 230, 231, 230, 230, 230, 230, 231, 231, 229, 230, 230, 231, 231, 230, 230, 230, 230, 230, 231, 230, 229, 230, 231, 231, 230, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 231, 230, 230, 232, 232, 232, 231, 231, 232, 232, 232, 232, 231, 231, 233, 232, 233, 232, 232, 232, 234, 234, 234, 234, 234, 235, 236, 236, 232, 227, 211, 161, 161, 157, 156, 158, 163, 159, 153, 151, 140, 144, 140, 144, 136, 150, 182, 187, 189, 166, 160, 175, 150, 82, 49, 46, 58, 79, 142, 167, 151, 59, 129, 166, 160, 98, 58, 117, 161, 166, 132, 156, 71, 42, 45, 68, 147, 146, 43, 42, 53, 135, 153, 101, 52, 52, 68, 129, 213, 231, 235, 236, 236, 234, 224, 187, 133, 54, 65, 50, 46, 56, 108, 209, 229, 229, 229, 229, 230, 231, 231, 230, 228, 229, 231, 232, 230, 230, 229, 230, 229, 230, 229, 229, 230, 231, 231, 229, 229, 228, 230, 230, 231, 229, 230, 229, 231, 231, 230, 229, 225, 222, 217, 224, 223, 219, 217, 125, 215, 224, 223, 221, 224, 220, 224, 224, 225, 226, 226, 225, 228, 227, 227, 227, 225, 228, 228, 228, 226, 227, 228, 228, 227, 227, 226, 226, 227, 228, 227, 226, 225, 227, 228, 228, 225, 226, 227, 229, 230, 230, 228, 229, 230, 231, 231, 229, 230, 229, 230, 230, 229, 229, 229, 229, 230, 230, 230, 230, 229, 231, 232, 231, 229, 230, 230, 231, 231, 230, 230, 229, 230, 230, 231, 229, 229, 229, 231, 230, 231, 230, 230, 230, 232, 231, 230, 229, 230, 231, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 230, 231, 230, 232, 231, 232, 231, 231, 231, 233, 233, 232, 232, 232, 233, 233, 233, 232, 233, 233, 234, 234, 234, 234, 234, 235, 236, 235, 231, 222, 175, 171, 165, 167, 160, 162, 162, 155, 149, 146, 139, 149, 140, 133, 137, 167, 192, 199, 185, 158, 175, 164, 105, 51, 38, 42, 50, 75, 129, 171, 157, 69, 106, 165, 158, 91, 76, 97, 167, 166, 78, 150, 105, 45, 48, 75, 146, 140, 44, 46, 56, 131, 165, 122, 42, 39, 48, 72, 120, 208, 232, 235, 236, 236, 232, 222, 181, 121, 52, 48, 47, 61, 137, 214, 227, 229, 229, 229, 230, 230, 231, 230, 229, 229, 231, 231, 230, 230, 230, 231, 231, 231, 229, 228, 229, 230, 231, 230, 228, 228, 229, 230, 231, 230, 230, 230, 231, 230, 230, 229, 224, 222, 218, 228, 223, 220, 219, 135, 213, 223, 223, 223, 224, 221, 224, 223, 225, 226, 224, 225, 225, 227, 226, 224, 224, 226, 226, 227, 227, 225, 226, 225, 226, 228, 227, 227, 227, 229, 227, 226, 227, 227, 228, 229, 228, 226, 227, 229, 230, 230, 229, 229, 229, 231, 231, 230, 229, 229, 230, 230, 229, 229, 228, 229, 229, 230, 230, 230, 229, 230, 231, 231, 229, 230, 230, 231, 231, 231, 229, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 229, 230, 230, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 232, 232, 232, 230, 231, 231, 232, 232, 232, 231, 231, 232, 233, 233, 232, 233, 233, 234, 234, 235, 234, 234, 235, 235, 233, 227, 180, 174, 169, 167, 162, 167, 165, 155, 152, 149, 146, 148, 144, 134, 134, 161, 187, 200, 198, 169, 171, 178, 133, 55, 52, 45, 46, 48, 83, 99, 177, 168, 88, 91, 166, 163, 64, 92, 88, 160, 163, 66, 91, 137, 87, 65, 101, 157, 99, 38, 39, 61, 110, 160, 126, 40, 34, 39, 47, 67, 112, 210, 232, 235, 236, 235, 231, 217, 168, 107, 50, 49, 59, 112, 189, 223, 228, 229, 229, 229, 230, 231, 230, 229, 229, 231, 231, 231, 230, 229, 230, 231, 231, 229, 228, 227, 230, 231, 230, 229, 228, 229, 230, 231, 230, 229, 229, 231, 229, 228, 230, 226, 223, 219, 228, 224, 225, 222, 119, 212, 224, 223, 223, 221, 221, 220, 224, 227, 225, 225, 226, 227, 226, 225, 224, 226, 226, 228, 228, 227, 225, 227, 228, 226, 227, 227, 227, 228, 230, 229, 228, 227, 226, 229, 228, 228, 228, 228, 229, 230, 230, 229, 230, 229, 231, 231, 230, 228, 229, 230, 230, 230, 229, 229, 229, 230, 230, 229, 229, 229, 230, 230, 231, 230, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 230, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 232, 231, 230, 230, 232, 232, 232, 231, 231, 231, 232, 232, 231, 232, 231, 232, 233, 232, 231, 232, 232, 233, 233, 233, 233, 233, 234, 234, 235, 234, 234, 235, 234, 230, 196, 176, 170, 169, 168, 166, 166, 162, 157, 149, 144, 150, 150, 130, 127, 145, 182, 193, 201, 187, 164, 185, 163, 81, 47, 46, 44, 47, 48, 60, 80, 174, 177, 87, 70, 160, 164, 68, 77, 111, 150, 156, 73, 51, 67, 82, 101, 139, 114, 48, 39, 41, 60, 97, 162, 135, 39, 34, 41, 38, 48, 72, 124, 217, 234, 235, 236, 234, 228, 209, 155, 79, 47, 50, 73, 140, 204, 224, 228, 228, 229, 231, 230, 230, 229, 230, 231, 231, 231, 229, 229, 229, 230, 231, 229, 229, 229, 229, 230, 231, 230, 228, 229, 231, 231, 231, 230, 229, 229, 230, 229, 228, 225, 223, 218, 228, 223, 224, 222, 126, 210, 221, 222, 223, 221, 223, 223, 225, 227, 224, 226, 225, 227, 226, 227, 226, 224, 226, 227, 227, 226, 227, 228, 226, 225, 226, 226, 226, 227, 229, 229, 226, 226, 228, 229, 228, 228, 228, 228, 229, 230, 229, 229, 229, 229, 230, 231, 230, 229, 229, 230, 231, 230, 229, 229, 229, 231, 230, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 232, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 231, 232, 232, 232, 233, 232, 231, 232, 233, 233, 233, 233, 233, 233, 235, 234, 235, 235, 234, 234, 231, 216, 177, 174, 173, 170, 176, 172, 171, 159, 149, 154, 152, 155, 154, 128, 136, 170, 193, 199, 201, 174, 179, 177, 119, 50, 46, 46, 44, 43, 44, 56, 68, 158, 172, 92, 62, 161, 164, 71, 64, 118, 141, 152, 82, 53, 73, 106, 97, 63, 48, 48, 41, 44, 50, 80, 158, 142, 44, 37, 38, 36, 39, 53, 72, 146, 225, 234, 236, 235, 232, 226, 194, 134, 57, 46, 56, 84, 160, 212, 226, 227, 227, 229, 231, 230, 230, 231, 231, 231, 230, 229, 229, 230, 231, 231, 230, 229, 229, 228, 230, 230, 230, 227, 230, 231, 232, 231, 229, 228, 230, 228, 228, 227, 225, 224, 219, 227, 224, 221, 222, 115, 212, 224, 221, 220, 221, 221, 225, 226, 226, 223, 227, 226, 227, 227, 226, 224, 224, 226, 228, 228, 227, 227, 228, 227, 226, 227, 228, 228, 228, 228, 229, 228, 227, 227, 229, 228, 229, 228, 228, 228, 229, 230, 229, 230, 230, 230, 231, 230, 229, 230, 230, 231, 230, 229, 229, 229, 231, 231, 230, 230, 230, 231, 231, 232, 230, 230, 230, 231, 231, 231, 229, 230, 230, 231, 230, 230, 230, 229, 231, 231, 230, 230, 230, 230, 231, 231, 230, 229, 229, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 232, 230, 230, 231, 232, 232, 231, 231, 230, 231, 232, 232, 231, 231, 231, 233, 233, 232, 231, 231, 233, 233, 233, 232, 233, 233, 235, 234, 235, 235, 233, 231, 227, 178, 183, 174, 173, 173, 175, 172, 166, 155, 155, 156, 165, 169, 160, 148, 154, 185, 200, 199, 189, 170, 186, 158, 64, 54, 43, 49, 48, 42, 48, 58, 66, 158, 170, 95, 64, 165, 165, 77, 58, 81, 155, 138, 86, 70, 117, 68, 46, 48, 41, 41, 39, 41, 51, 68, 156, 144, 63, 36, 35, 38, 35, 41, 57, 80, 180, 231, 235, 235, 234, 232, 223, 174, 105, 46, 55, 61, 108, 188, 220, 228, 227, 229, 230, 230, 230, 231, 231, 231, 230, 229, 229, 231, 230, 231, 230, 229, 229, 230, 230, 230, 230, 228, 230, 231, 230, 229, 227, 229, 230, 230, 227, 228, 223, 220, 216, 227, 222, 220, 224, 122, 214, 226, 224, 221, 222, 221, 226, 227, 226, 223, 225, 225, 226, 227, 224, 226, 224, 228, 228, 227, 228, 227, 228, 228, 229, 228, 228, 227, 229, 229, 229, 228, 226, 228, 230, 229, 228, 228, 226, 227, 229, 229, 230, 229, 229, 230, 230, 230, 229, 229, 231, 230, 230, 229, 228, 229, 231, 231, 230, 230, 230, 231, 230, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 232, 231, 230, 230, 232, 232, 232, 231, 231, 231, 233, 233, 232, 231, 231, 232, 233, 233, 233, 233, 233, 234, 234, 235, 234, 232, 229, 195, 181, 179, 177, 174, 176, 176, 167, 161, 158, 158, 170, 170, 170, 178, 161, 173, 194, 199, 199, 173, 178, 178, 113, 48, 47, 49, 47, 52, 43, 46, 56, 61, 162, 174, 89, 74, 156, 164, 77, 56, 64, 155, 130, 88, 136, 145, 132, 106, 103, 89, 95, 52, 45, 48, 62, 159, 148, 58, 39, 39, 38, 38, 40, 56, 61, 88, 200, 233, 235, 235, 235, 229, 209, 148, 64, 46, 52, 72, 141, 203, 221, 226, 228, 230, 230, 230, 231, 231, 230, 230, 229, 229, 230, 230, 231, 230, 230, 230, 230, 231, 229, 229, 229, 230, 231, 230, 230, 229, 228, 229, 229, 229, 228, 224, 222, 215, 229, 223, 220, 224, 124, 216, 226, 226, 223, 222, 223, 225, 228, 226, 225, 227, 227, 224, 227, 225, 226, 227, 228, 230, 228, 228, 227, 226, 228, 227, 228, 228, 228, 229, 228, 228, 229, 228, 228, 230, 229, 227, 228, 228, 227, 229, 229, 230, 229, 229, 230, 231, 229, 229, 229, 230, 231, 229, 229, 229, 229, 231, 231, 230, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 229, 230, 231, 231, 231, 229, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 229, 229, 230, 230, 230, 231, 229, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 232, 230, 230, 230, 232, 232, 232, 231, 231, 232, 233, 233, 232, 232, 232, 233, 234, 233, 232, 233, 233, 234, 235, 235, 233, 229, 221, 173, 179, 178, 176, 181, 181, 179, 169, 162, 158, 167, 174, 179, 176, 175, 181, 188, 196, 202, 191, 167, 183, 165, 70, 50, 51, 57, 46, 45, 41, 42, 51, 54, 147, 168, 105, 63, 156, 162, 87, 56, 59, 149, 147, 112, 132, 166, 174, 165, 162, 166, 151, 55, 43, 50, 58, 162, 154, 63, 35, 37, 34, 36, 40, 38, 46, 67, 121, 221, 235, 235, 236, 233, 225, 184, 115, 50, 47, 58, 88, 170, 212, 224, 227, 230, 230, 230, 230, 232, 230, 230, 229, 230, 230, 231, 231, 229, 230, 230, 231, 230, 229, 229, 229, 230, 231, 230, 229, 230, 229, 230, 230, 231, 229, 225, 222, 214, 226, 222, 221, 226, 125, 218, 225, 226, 222, 222, 224, 226, 227, 228, 226, 226, 226, 226, 227, 226, 226, 228, 228, 230, 228, 228, 227, 227, 227, 227, 226, 227, 228, 230, 229, 229, 228, 228, 229, 229, 230, 229, 229, 227, 228, 230, 230, 229, 230, 229, 230, 231, 229, 229, 229, 230, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 230, 231, 230, 230, 229, 231, 231, 231, 229, 230, 230, 231, 232, 230, 230, 230, 230, 231, 231, 230, 229, 229, 231, 231, 231, 230, 230, 230, 231, 232, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 231, 231, 230, 230, 232, 231, 232, 231, 231, 232, 233, 233, 232, 232, 232, 233, 233, 234, 233, 233, 233, 235, 236, 234, 232, 229, 186, 180, 180, 179, 174, 175, 178, 172, 168, 162, 159, 172, 176, 179, 178, 180, 181, 187, 198, 203, 180, 176, 177, 140, 85, 80, 130, 131, 62, 43, 47, 42, 51, 55, 144, 172, 113, 59, 153, 173, 104, 54, 55, 142, 125, 97, 101, 128, 141, 143, 149, 142, 100, 49, 41, 50, 58, 152, 160, 58, 36, 39, 41, 43, 47, 41, 46, 59, 85, 173, 230, 235, 236, 236, 230, 212, 155, 73, 45, 49, 67, 123, 189, 219, 225, 230, 230, 230, 230, 231, 230, 229, 229, 229, 230, 230, 230, 230, 229, 230, 231, 231, 230, 229, 229, 230, 231, 230, 228, 229, 228, 229, 229, 229, 230, 225, 223, 218, 225, 222, 220, 224, 114, 217, 225, 227, 224, 223, 225, 227, 227, 226, 226, 227, 226, 227, 228, 228, 226, 228, 228, 229, 228, 229, 227, 228, 228, 227, 227, 227, 227, 230, 229, 229, 228, 229, 229, 230, 230, 229, 229, 228, 228, 230, 230, 229, 230, 230, 231, 231, 230, 229, 229, 230, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 229, 229, 229, 231, 231, 231, 229, 230, 230, 232, 232, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 230, 230, 232, 232, 232, 231, 231, 232, 233, 233, 232, 232, 232, 233, 233, 233, 232, 233, 234, 235, 235, 233, 229, 218, 172, 180, 180, 176, 171, 180, 175, 171, 165, 157, 167, 179, 180, 182, 179, 178, 182, 193, 201, 195, 174, 184, 180, 104, 170, 103, 169, 168, 75, 48, 48, 42, 52, 55, 141, 170, 131, 62, 140, 180, 134, 54, 57, 90, 56, 54, 71, 81, 57, 53, 64, 78, 46, 38, 37, 50, 52, 153, 165, 67, 42, 60, 126, 94, 90, 115, 70, 54, 83, 125, 212, 234, 236, 236, 234, 226, 182, 126, 51, 49, 57, 80, 160, 213, 225, 229, 230, 230, 230, 230, 230, 230, 229, 229, 229, 230, 231, 229, 228, 230, 229, 230, 230, 228, 228, 229, 231, 228, 229, 229, 229, 230, 230, 229, 229, 226, 225, 221, 228, 222, 222, 223, 114, 218, 227, 226, 223, 225, 226, 225, 227, 228, 225, 228, 227, 229, 227, 228, 228, 229, 229, 229, 229, 228, 227, 229, 230, 228, 228, 227, 228, 230, 229, 229, 229, 229, 230, 230, 230, 229, 228, 229, 229, 230, 231, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 231, 230, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 230, 230, 229, 230, 231, 231, 230, 230, 229, 231, 232, 231, 230, 230, 230, 232, 232, 231, 230, 230, 231, 232, 232, 231, 230, 230, 232, 233, 232, 231, 232, 232, 232, 233, 232, 232, 232, 233, 233, 233, 232, 233, 234, 236, 234, 232, 227, 184, 174, 179, 178, 177, 175, 179, 175, 172, 161, 163, 178, 180, 180, 180, 184, 184, 190, 199, 202, 196, 167, 186, 159, 71, 88, 103, 161, 170, 83, 48, 77, 68, 66, 57, 112, 137, 111, 56, 113, 152, 125, 54, 66, 100, 48, 48, 68, 91, 93, 50, 51, 82, 60, 41, 45, 67, 67, 136, 158, 73, 46, 118, 139, 48, 51, 105, 151, 77, 98, 192, 158, 230, 235, 236, 236, 229, 213, 159, 76, 49, 52, 63, 119, 196, 223, 229, 229, 230, 229, 230, 231, 230, 229, 228, 229, 230, 230, 229, 228, 229, 230, 230, 229, 229, 229, 231, 230, 231, 230, 230, 229, 230, 230, 230, 228, 226, 226, 220, 229, 223, 220, 222, 129, 216, 228, 228, 225, 225, 228, 227, 226, 225, 226, 226, 227, 230, 227, 228, 228, 228, 229, 229, 228, 227, 226, 229, 229, 229, 229, 228, 228, 229, 229, 229, 229, 229, 229, 231, 231, 230, 228, 229, 229, 230, 230, 229, 230, 229, 230, 230, 229, 230, 230, 231, 231, 231, 230, 230, 230, 231, 230, 230, 229, 229, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 230, 229, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 230, 232, 232, 230, 230, 230, 232, 231, 231, 231, 230, 231, 232, 232, 231, 231, 230, 231, 232, 232, 232, 232, 232, 233, 233, 233, 232, 232, 233, 234, 233, 233, 233, 234, 235, 233, 229, 223, 164, 177, 180, 181, 173, 179, 175, 169, 171, 165, 173, 180, 182, 181, 182, 184, 188, 189, 202, 206, 191, 177, 182, 149, 63, 59, 90, 160, 174, 99, 108, 128, 58, 120, 92, 57, 47, 51, 48, 46, 54, 55, 58, 90, 135, 52, 50, 100, 98, 96, 71, 63, 131, 122, 39, 44, 60, 70, 54, 61, 46, 46, 144, 131, 46, 50, 72, 151, 117, 57, 87, 97, 208, 235, 236, 236, 232, 225, 186, 115, 50, 47, 57, 85, 172, 219, 229, 230, 229, 230, 231, 231, 230, 229, 229, 230, 230, 230, 229, 229, 230, 230, 231, 229, 230, 229, 230, 231, 231, 230, 229, 230, 230, 230, 229, 228, 225, 224, 222, 225, 222, 217, 221, 121, 216, 226, 226, 225, 226, 226, 228, 226, 226, 226, 227, 228, 229, 229, 228, 228, 227, 229, 228, 228, 228, 228, 229, 229, 229, 229, 229, 227, 229, 229, 229, 229, 229, 229, 230, 231, 229, 229, 229, 229, 230, 231, 230, 229, 230, 230, 230, 230, 230, 229, 230, 230, 230, 230, 230, 229, 231, 231, 230, 229, 229, 231, 230, 230, 229, 229, 230, 231, 231, 231, 230, 229, 230, 231, 230, 230, 229, 230, 231, 231, 230, 229, 229, 230, 231, 230, 229, 229, 229, 230, 231, 230, 230, 230, 230, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 232, 233, 233, 232, 232, 232, 232, 234, 233, 233, 233, 234, 235, 233, 228, 201, 178, 175, 183, 180, 176, 176, 174, 169, 173, 168, 178, 184, 183, 186, 186, 185, 187, 193, 205, 207, 182, 180, 176, 121, 53, 59, 59, 152, 182, 108, 153, 120, 61, 101, 152, 63, 47, 47, 45, 42, 42, 48, 49, 51, 94, 50, 47, 51, 58, 54, 61, 82, 75, 62, 42, 45, 46, 48, 99, 93, 43, 42, 137, 143, 48, 51, 73, 142, 135, 46, 59, 83, 161, 232, 236, 237, 234, 228, 209, 150, 61, 48, 50, 69, 137, 207, 227, 229, 230, 230, 231, 231, 230, 230, 230, 230, 231, 230, 229, 229, 230, 230, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 230, 230, 228, 230, 225, 225, 221, 228, 222, 219, 223, 123, 218, 226, 226, 224, 226, 226, 228, 227, 226, 226, 226, 227, 229, 229, 228, 228, 227, 228, 228, 229, 229, 228, 230, 230, 229, 229, 228, 229, 230, 230, 230, 229, 229, 229, 230, 230, 230, 230, 230, 230, 230, 231, 230, 230, 230, 230, 231, 230, 230, 229, 231, 231, 230, 230, 230, 230, 231, 231, 229, 228, 229, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 229, 230, 231, 231, 231, 230, 230, 229, 230, 231, 230, 230, 230, 230, 231, 231, 229, 229, 230, 231, 231, 231, 230, 230, 231, 232, 231, 231, 231, 231, 232, 232, 232, 232, 232, 232, 233, 233, 232, 232, 232, 233, 234, 234, 233, 234, 235, 234, 232, 229, 175, 177, 176, 182, 178, 179, 178, 173, 175, 172, 171, 178, 181, 186, 186, 187, 187, 188, 200, 207, 205, 180, 190, 172, 110, 53, 53, 59, 141, 182, 123, 164, 112, 66, 84, 162, 99, 51, 46, 46, 39, 43, 44, 48, 57, 109, 110, 49, 48, 43, 47, 52, 57, 138, 78, 41, 42, 43, 38, 38, 39, 41, 48, 96, 150, 91, 62, 72, 148, 110, 49, 51, 76, 106, 218, 236, 236, 235, 230, 222, 178, 82, 48, 44, 63, 95, 192, 224, 229, 230, 230, 231, 231, 230, 230, 229, 230, 230, 231, 229, 230, 230, 230, 230, 230, 230, 229, 230, 231, 230, 230, 229, 229, 231, 230, 229, 229, 226, 225, 218, 229, 224, 223, 223, 125, 217, 225, 226, 224, 226, 226, 228, 228, 227, 227, 227, 228, 229, 229, 229, 229, 228, 229, 228, 229, 228, 227, 229, 230, 230, 230, 229, 230, 230, 230, 230, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 229, 229, 231, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 229, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 230, 231, 231, 232, 232, 232, 231, 232, 232, 233, 232, 232, 231, 233, 234, 234, 233, 234, 234, 233, 229, 218, 171, 178, 178, 182, 178, 178, 178, 174, 175, 177, 179, 180, 187, 183, 190, 189, 189, 196, 205, 203, 206, 182, 184, 167, 79, 48, 53, 57, 136, 184, 137, 166, 122, 63, 70, 162, 124, 50, 43, 43, 43, 45, 50, 51, 47, 89, 93, 59, 50, 51, 53, 59, 67, 121, 104, 57, 45, 41, 41, 39, 39, 43, 46, 51, 95, 123, 96, 109, 124, 56, 48, 50, 66, 84, 183, 234, 236, 235, 233, 227, 200, 122, 49, 44, 52, 78, 168, 219, 229, 230, 230, 230, 231, 230, 230, 230, 230, 230, 230, 229, 230, 230, 231, 231, 231, 230, 229, 230, 230, 230, 230, 230, 229, 229, 230, 230, 230, 227, 225, 221, 229, 225, 223, 224, 129, 219, 226, 227, 224, 224, 225, 226, 225, 226, 226, 228, 228, 230, 230, 229, 228, 227, 228, 230, 229, 229, 228, 229, 231, 230, 230, 230, 229, 230, 230, 230, 229, 230, 230, 232, 231, 230, 230, 229, 231, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 230, 230, 230, 229, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 229, 229, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 231, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 233, 231, 231, 231, 232, 233, 233, 231, 232, 233, 234, 234, 233, 234, 233, 233, 229, 193, 177, 178, 182, 182, 180, 183, 185, 177, 178, 175, 180, 182, 188, 187, 188, 193, 192, 196, 204, 207, 205, 178, 186, 159, 59, 52, 52, 60, 124, 183, 145, 155, 139, 62, 66, 151, 129, 52, 49, 45, 45, 45, 43, 43, 49, 48, 78, 128, 79, 61, 72, 84, 110, 69, 55, 64, 62, 48, 41, 42, 45, 40, 44, 46, 50, 77, 102, 85, 54, 50, 48, 48, 61, 81, 132, 229, 235, 235, 234, 228, 216, 151, 57, 44, 48, 68, 132, 207, 228, 229, 230, 231, 231, 230, 230, 229, 230, 230, 230, 230, 230, 230, 231, 231, 230, 230, 230, 230, 230, 231, 229, 230, 229, 228, 229, 230, 230, 228, 227, 221, 226, 224, 223, 224, 140, 219, 228, 225, 226, 225, 227, 226, 227, 227, 227, 228, 227, 229, 230, 229, 227, 227, 229, 230, 229, 228, 229, 229, 230, 230, 230, 229, 228, 231, 230, 230, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 230, 230, 229, 229, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 229, 230, 229, 231, 231, 231, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 232, 231, 231, 231, 232, 232, 233, 232, 231, 232, 232, 233, 233, 232, 232, 233, 234, 234, 233, 234, 233, 232, 229, 179, 178, 175, 186, 181, 178, 186, 182, 175, 178, 181, 182, 184, 183, 189, 189, 193, 195, 197, 207, 209, 200, 181, 187, 148, 55, 50, 51, 61, 122, 177, 149, 134, 152, 65, 67, 159, 100, 48, 46, 41, 40, 41, 42, 46, 43, 49, 48, 102, 90, 128, 130, 83, 91, 46, 50, 49, 60, 57, 49, 40, 40, 44, 42, 48, 95, 87, 62, 57, 56, 67, 52, 49, 57, 74, 104, 216, 235, 235, 235, 231, 224, 176, 82, 44, 45, 75, 94, 191, 224, 229, 230, 230, 231, 230, 229, 229, 230, 230, 230, 230, 229, 230, 231, 231, 231, 229, 229, 230, 231, 231, 229, 229, 229, 229, 230, 230, 229, 227, 226, 220, 225, 222, 222, 224, 135, 220, 228, 228, 226, 225, 226, 224, 226, 227, 228, 227, 229, 229, 230, 227, 229, 228, 228, 229, 228, 229, 229, 228, 229, 230, 230, 229, 229, 231, 231, 230, 229, 230, 230, 231, 231, 230, 230, 229, 230, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 232, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 232, 231, 231, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 232, 231, 231, 231, 231, 232, 232, 232, 231, 232, 233, 233, 232, 232, 232, 234, 234, 234, 234, 233, 233, 229, 220, 168, 175, 179, 188, 177, 188, 185, 182, 180, 179, 183, 185, 184, 181, 187, 189, 194, 196, 202, 206, 210, 201, 181, 181, 137, 48, 49, 52, 64, 106, 176, 159, 74, 152, 91, 84, 146, 59, 41, 44, 41, 42, 39, 41, 41, 46, 47, 50, 51, 93, 78, 67, 71, 61, 51, 45, 42, 51, 43, 56, 46, 37, 49, 46, 64, 158, 162, 161, 155, 153, 123, 50, 55, 58, 72, 95, 188, 234, 235, 235, 233, 227, 191, 111, 50, 48, 56, 83, 176, 222, 230, 230, 231, 231, 231, 229, 230, 229, 231, 231, 229, 229, 230, 231, 230, 230, 230, 230, 230, 228, 230, 229, 229, 227, 230, 230, 231, 229, 228, 225, 222, 226, 224, 224, 224, 144, 219, 228, 227, 226, 226, 226, 227, 228, 228, 229, 229, 229, 230, 230, 228, 227, 227, 228, 230, 228, 228, 228, 228, 229, 230, 229, 229, 229, 231, 231, 230, 229, 229, 230, 231, 231, 230, 230, 229, 232, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 230, 229, 230, 231, 231, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 231, 230, 230, 230, 231, 231, 231, 229, 230, 231, 232, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 231, 231, 231, 231, 231, 233, 232, 231, 231, 232, 233, 233, 233, 232, 232, 233, 234, 234, 234, 233, 232, 228, 208, 175, 180, 180, 187, 181, 184, 187, 182, 184, 184, 184, 187, 184, 184, 193, 189, 195, 192, 202, 209, 214, 199, 186, 187, 138, 52, 48, 55, 58, 74, 125, 111, 56, 67, 87, 89, 67, 47, 43, 43, 37, 45, 39, 40, 39, 36, 44, 56, 92, 179, 161, 157, 174, 159, 99, 43, 47, 45, 41, 45, 54, 49, 46, 55, 80, 154, 163, 157, 157, 144, 87, 56, 55, 62, 69, 90, 148, 232, 235, 236, 234, 228, 203, 136, 52, 50, 56, 73, 145, 215, 228, 229, 231, 230, 230, 229, 229, 229, 230, 230, 229, 230, 228, 230, 231, 230, 230, 229, 229, 230, 230, 228, 227, 229, 231, 229, 229, 228, 228, 226, 220, 228, 221, 220, 223, 130, 218, 228, 227, 224, 226, 226, 227, 229, 228, 228, 229, 230, 230, 230, 228, 227, 227, 229, 230, 229, 228, 229, 229, 230, 230, 229, 229, 229, 230, 231, 230, 228, 229, 230, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 229, 229, 230, 230, 231, 231, 229, 230, 229, 231, 231, 230, 230, 229, 231, 231, 231, 229, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 232, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 232, 230, 230, 231, 232, 233, 232, 231, 231, 232, 233, 233, 233, 232, 232, 234, 234, 234, 234, 233, 232, 230, 191, 178, 179, 184, 186, 185, 187, 187, 182, 180, 180, 187, 184, 188, 189, 196, 192, 192, 193, 203, 210, 211, 199, 196, 189, 138, 55, 49, 49, 54, 50, 54, 52, 47, 51, 45, 47, 40, 40, 39, 41, 41, 56, 40, 40, 37, 40, 50, 56, 169, 170, 176, 180, 179, 150, 108, 49, 55, 52, 46, 53, 53, 53, 61, 53, 51, 61, 66, 56, 59, 57, 49, 55, 56, 61, 68, 90, 120, 223, 235, 235, 235, 229, 208, 150, 56, 52, 54, 68, 116, 206, 228, 229, 231, 231, 230, 229, 229, 230, 230, 229, 228, 229, 230, 231, 231, 231, 230, 229, 229, 230, 230, 229, 228, 229, 231, 231, 230, 229, 225, 225, 217, 228, 224, 221, 223, 146, 222, 227, 227, 226, 226, 226, 227, 227, 227, 226, 227, 229, 230, 230, 228, 228, 229, 229, 230, 229, 228, 229, 230, 230, 230, 230, 229, 230, 230, 231, 230, 229, 229, 230, 231, 231, 229, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 231, 232, 232, 230, 231, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 233, 232, 231, 231, 232, 233, 233, 232, 232, 232, 234, 234, 234, 234, 233, 231, 230, 189, 183, 183, 184, 188, 182, 191, 185, 177, 176, 182, 186, 191, 189, 188, 196, 192, 192, 193, 199, 208, 210, 196, 189, 185, 133, 46, 48, 53, 64, 89, 92, 89, 65, 49, 45, 44, 44, 43, 44, 39, 39, 38, 41, 39, 35, 41, 47, 61, 148, 166, 152, 137, 130, 100, 98, 52, 47, 50, 45, 47, 46, 53, 57, 63, 67, 49, 53, 47, 54, 50, 61, 64, 64, 66, 69, 84, 100, 212, 234, 235, 235, 230, 217, 159, 69, 51, 59, 69, 103, 199, 225, 229, 231, 231, 230, 230, 229, 230, 230, 231, 229, 230, 230, 231, 232, 231, 230, 229, 228, 230, 230, 229, 229, 230, 231, 231, 231, 230, 228, 225, 217, 228, 225, 220, 223, 127, 220, 228, 227, 227, 227, 228, 228, 229, 229, 228, 228, 228, 230, 230, 229, 229, 230, 230, 229, 228, 228, 229, 229, 230, 230, 230, 229, 230, 231, 231, 230, 229, 229, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 229, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 229, 229, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 233, 232, 231, 232, 232, 233, 233, 232, 232, 232, 233, 234, 234, 233, 233, 230, 230, 183, 180, 180, 186, 186, 185, 188, 183, 179, 179, 179, 186, 186, 188, 186, 192, 193, 190, 196, 202, 210, 211, 196, 189, 189, 135, 52, 53, 70, 142, 125, 89, 123, 146, 90, 51, 40, 40, 45, 43, 44, 39, 38, 44, 41, 41, 40, 48, 52, 124, 133, 126, 139, 169, 159, 131, 57, 47, 49, 46, 61, 48, 51, 47, 58, 59, 72, 67, 58, 60, 114, 142, 149, 143, 107, 68, 81, 104, 191, 233, 235, 235, 231, 221, 168, 82, 50, 52, 65, 96, 186, 224, 229, 231, 231, 230, 230, 229, 231, 230, 231, 230, 230, 230, 231, 230, 231, 229, 228, 230, 230, 230, 229, 229, 230, 231, 231, 231, 228, 228, 226, 219, 228, 224, 222, 224, 123, 217, 227, 228, 227, 227, 228, 227, 228, 229, 228, 226, 229, 230, 231, 228, 227, 228, 229, 229, 229, 228, 229, 229, 230, 230, 230, 229, 229, 231, 230, 231, 230, 229, 229, 231, 230, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 230, 231, 230, 229, 230, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 230, 230, 231, 231, 231, 231, 230, 230, 231, 232, 232, 231, 230, 231, 232, 232, 232, 231, 231, 232, 233, 232, 232, 232, 232, 233, 234, 234, 233, 233, 230, 230, 181, 181, 179, 185, 185, 184, 189, 184, 177, 179, 179, 186, 185, 185, 190, 185, 194, 192, 189, 198, 209, 211, 195, 191, 188, 142, 55, 59, 126, 165, 70, 57, 87, 140, 159, 61, 47, 46, 42, 43, 45, 38, 39, 43, 42, 44, 37, 44, 49, 54, 60, 101, 162, 173, 178, 159, 115, 56, 55, 50, 56, 56, 60, 55, 60, 65, 69, 110, 118, 81, 146, 163, 148, 163, 111, 106, 113, 127, 178, 231, 234, 234, 231, 224, 176, 90, 56, 56, 65, 90, 173, 222, 230, 231, 231, 231, 230, 230, 230, 229, 231, 230, 229, 230, 232, 231, 231, 229, 229, 230, 230, 230, 229, 229, 230, 231, 231, 230, 229, 228, 227, 219, 226, 224, 223, 223, 129, 219, 226, 227, 227, 227, 228, 229, 229, 228, 227, 228, 229, 229, 229, 226, 228, 227, 228, 229, 230, 228, 229, 230, 231, 231, 230, 229, 228, 230, 231, 230, 230, 229, 230, 231, 230, 230, 229, 229, 231, 231, 231, 229, 229, 230, 231, 231, 230, 229, 229, 230, 231, 230, 229, 230, 230, 230, 230, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 230, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 229, 230, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 232, 231, 230, 231, 232, 232, 232, 231, 231, 231, 233, 233, 232, 232, 233, 233, 234, 234, 232, 232, 230, 229, 179, 183, 182, 186, 186, 191, 190, 184, 180, 178, 179, 184, 183, 185, 187, 187, 188, 185, 188, 200, 206, 209, 199, 187, 188, 143, 56, 54, 141, 159, 59, 56, 65, 107, 166, 117, 43, 40, 39, 37, 40, 39, 37, 38, 40, 38, 40, 38, 44, 48, 57, 142, 166, 164, 163, 170, 161, 140, 143, 140, 142, 144, 148, 148, 143, 152, 153, 163, 174, 156, 150, 168, 194, 205, 200, 201, 204, 207, 210, 216, 231, 234, 232, 227, 180, 112, 57, 58, 66, 88, 166, 218, 229, 231, 231, 230, 230, 228, 230, 230, 230, 230, 230, 230, 232, 231, 230, 230, 229, 229, 228, 230, 227, 228, 229, 230, 231, 230, 230, 227, 226, 218, 227, 223, 221, 224, 118, 218, 227, 226, 225, 227, 228, 228, 228, 228, 227, 228, 228, 229, 229, 228, 228, 227, 229, 229, 229, 229, 229, 230, 230, 231, 230, 229, 228, 230, 231, 230, 229, 229, 229, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 229, 229, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 231, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 232, 232, 231, 230, 231, 231, 232, 232, 231, 232, 231, 233, 233, 233, 232, 232, 233, 234, 234, 233, 232, 230, 230, 185, 181, 182, 187, 186, 189, 192, 183, 179, 178, 179, 185, 187, 184, 183, 183, 189, 190, 188, 201, 207, 211, 203, 182, 191, 155, 61, 54, 126, 155, 72, 53, 58, 86, 161, 154, 51, 38, 40, 40, 40, 42, 41, 33, 37, 35, 39, 38, 45, 70, 68, 145, 165, 166, 140, 174, 170, 171, 169, 166, 167, 158, 158, 152, 150, 151, 146, 144, 145, 146, 128, 143, 160, 160, 168, 146, 134, 148, 158, 222, 232, 234, 233, 228, 182, 122, 59, 55, 66, 88, 154, 217, 229, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 231, 231, 230, 231, 229, 229, 230, 228, 228, 229, 228, 228, 230, 230, 230, 229, 229, 226, 220, 228, 224, 222, 224, 112, 215, 226, 218, 227, 227, 227, 228, 228, 229, 228, 228, 229, 229, 228, 227, 228, 227, 230, 229, 229, 229, 227, 229, 229, 231, 230, 229, 229, 230, 230, 230, 229, 230, 229, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 229, 230, 230, 231, 230, 229, 229, 231, 231, 231, 230, 230, 230, 232, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 231, 231, 232, 233, 232, 231, 232, 233, 233, 232, 232, 232, 233, 234, 234, 234, 232, 230, 230, 186, 183, 185, 188, 181, 186, 193, 181, 183, 179, 179, 181, 182, 182, 185, 186, 189, 189, 191, 197, 209, 217, 208, 189, 197, 166, 78, 54, 78, 152, 118, 61, 61, 76, 160, 161, 51, 43, 43, 40, 40, 42, 37, 45, 42, 39, 39, 37, 47, 53, 59, 150, 174, 176, 163, 169, 163, 120, 99, 93, 90, 85, 79, 67, 68, 62, 61, 59, 63, 83, 101, 110, 96, 92, 140, 144, 90, 144, 168, 225, 234, 234, 232, 226, 185, 119, 61, 61, 68, 100, 147, 215, 228, 230, 231, 230, 229, 229, 230, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 229, 229, 230, 229, 229, 228, 230, 230, 230, 230, 230, 226, 220, 227, 224, 224, 223, 146, 217, 227, 224, 225, 225, 225, 227, 228, 230, 227, 228, 228, 229, 227, 228, 228, 228, 229, 230, 230, 229, 228, 228, 230, 230, 231, 230, 230, 230, 231, 230, 229, 229, 229, 231, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 231, 230, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 232, 230, 231, 232, 232, 233, 232, 232, 231, 233, 233, 233, 232, 232, 233, 234, 234, 234, 232, 231, 230, 185, 182, 184, 186, 182, 184, 186, 182, 182, 182, 180, 183, 184, 184, 187, 186, 187, 190, 194, 199, 212, 218, 213, 187, 195, 168, 68, 44, 55, 86, 124, 96, 76, 63, 159, 156, 51, 42, 42, 44, 43, 43, 43, 41, 41, 41, 41, 39, 44, 49, 59, 96, 161, 170, 170, 166, 134, 59, 50, 48, 49, 54, 56, 51, 52, 50, 52, 55, 57, 105, 94, 57, 67, 72, 99, 137, 95, 98, 115, 222, 233, 234, 232, 227, 189, 124, 63, 57, 69, 95, 148, 211, 229, 231, 231, 231, 230, 229, 230, 230, 230, 230, 230, 230, 231, 231, 231, 229, 229, 228, 229, 230, 229, 228, 228, 229, 230, 230, 229, 229, 226, 220, 226, 225, 224, 224, 134, 216, 228, 227, 225, 225, 227, 227, 229, 230, 227, 227, 227, 228, 229, 226, 227, 226, 229, 230, 230, 228, 229, 228, 230, 231, 231, 230, 229, 230, 231, 231, 230, 229, 229, 231, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 231, 230, 230, 229, 230, 230, 231, 231, 230, 230, 229, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 231, 229, 230, 231, 231, 231, 230, 230, 230, 231, 232, 230, 230, 230, 231, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 232, 232, 233, 233, 233, 232, 232, 234, 235, 234, 234, 233, 231, 230, 185, 177, 179, 189, 181, 182, 193, 182, 179, 179, 183, 182, 184, 184, 187, 188, 185, 190, 194, 200, 211, 222, 216, 192, 199, 179, 90, 49, 54, 103, 113, 58, 58, 79, 163, 111, 43, 39, 44, 43, 43, 43, 42, 57, 42, 39, 40, 40, 47, 56, 68, 57, 106, 146, 157, 156, 74, 54, 49, 49, 48, 49, 51, 48, 49, 50, 53, 55, 59, 96, 95, 55, 57, 67, 107, 158, 112, 120, 119, 220, 233, 234, 232, 224, 179, 119, 58, 66, 68, 97, 152, 217, 229, 231, 231, 230, 230, 229, 230, 231, 230, 231, 229, 230, 231, 231, 231, 230, 230, 229, 230, 230, 229, 228, 228, 229, 230, 231, 229, 229, 226, 220, 227, 224, 223, 225, 125, 217, 226, 225, 224, 225, 226, 226, 227, 229, 226, 226, 226, 228, 228, 226, 226, 227, 229, 230, 230, 229, 228, 229, 230, 231, 230, 229, 230, 230, 230, 230, 230, 229, 230, 230, 231, 231, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 229, 230, 230, 232, 231, 230, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 229, 229, 231, 230, 231, 230, 230, 230, 231, 230, 229, 229, 229, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 232, 233, 233, 233, 232, 232, 234, 234, 234, 233, 233, 231, 230, 195, 178, 181, 186, 185, 187, 192, 184, 178, 178, 177, 182, 184, 184, 186, 186, 192, 194, 194, 204, 212, 222, 216, 194, 196, 183, 100, 50, 52, 112, 148, 79, 64, 134, 144, 55, 45, 45, 43, 42, 38, 41, 43, 45, 45, 44, 41, 40, 44, 46, 47, 46, 59, 70, 128, 158, 106, 54, 43, 51, 50, 50, 49, 45, 51, 52, 54, 54, 58, 65, 108, 75, 61, 71, 138, 146, 76, 99, 122, 204, 230, 233, 231, 224, 179, 116, 61, 63, 77, 108, 156, 217, 229, 231, 232, 231, 229, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 230, 229, 228, 229, 230, 230, 230, 230, 226, 229, 225, 220, 227, 225, 223, 224, 130, 220, 224, 226, 224, 224, 225, 226, 227, 228, 226, 226, 227, 228, 228, 227, 228, 228, 227, 230, 228, 228, 228, 229, 230, 231, 229, 229, 230, 231, 230, 231, 230, 229, 229, 230, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 229, 230, 230, 232, 231, 231, 229, 229, 230, 230, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 232, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 231, 232, 230, 234, 231, 231, 231, 230, 231, 231, 231, 231, 230, 230, 232, 232, 231, 230, 230, 231, 231, 231, 231, 230, 231, 232, 232, 231, 231, 231, 232, 233, 233, 233, 232, 232, 233, 234, 234, 233, 233, 231, 230, 191, 179, 181, 189, 187, 185, 191, 185, 181, 179, 181, 182, 181, 189, 187, 189, 192, 194, 196, 202, 210, 221, 222, 197, 196, 204, 127, 49, 47, 53, 99, 110, 110, 118, 57, 43, 44, 41, 39, 40, 40, 40, 43, 44, 47, 40, 46, 39, 41, 47, 42, 47, 50, 63, 88, 163, 147, 58, 50, 47, 51, 47, 49, 49, 46, 50, 49, 58, 56, 60, 69, 103, 96, 111, 124, 82, 74, 86, 112, 221, 232, 230, 227, 217, 175, 111, 67, 65, 79, 116, 163, 217, 230, 230, 231, 231, 230, 229, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 230, 229, 230, 230, 228, 229, 229, 230, 228, 228, 227, 225, 219, 226, 223, 221, 225, 124, 220, 225, 228, 225, 225, 226, 227, 229, 229, 226, 225, 227, 228, 228, 227, 227, 227, 228, 230, 230, 229, 229, 230, 230, 230, 229, 229, 229, 231, 231, 230, 229, 229, 229, 230, 230, 229, 228, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 229, 230, 230, 231, 230, 230, 230, 231, 231, 230, 230, 229, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 232, 231, 230, 230, 232, 232, 231, 230, 230, 230, 231, 230, 231, 230, 230, 231, 232, 231, 230, 230, 230, 232, 232, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 231, 231, 231, 231, 231, 232, 232, 231, 231, 232, 233, 233, 232, 232, 233, 232, 234, 234, 233, 233, 232, 231, 203, 184, 184, 192, 191, 188, 192, 186, 182, 179, 179, 183, 187, 185, 188, 190, 193, 192, 193, 200, 212, 218, 224, 205, 194, 220, 164, 53, 46, 45, 47, 49, 47, 46, 43, 41, 42, 48, 41, 47, 42, 41, 43, 40, 46, 43, 42, 43, 40, 41, 45, 58, 48, 92, 66, 138, 161, 105, 49, 58, 52, 49, 48, 49, 53, 51, 51, 53, 50, 50, 53, 61, 58, 62, 63, 58, 69, 94, 117, 224, 234, 233, 229, 217, 172, 109, 67, 68, 83, 122, 164, 218, 230, 231, 231, 231, 230, 230, 231, 231, 230, 230, 230, 230, 232, 231, 230, 230, 229, 230, 230, 230, 230, 226, 228, 230, 231, 229, 228, 227, 226, 221, 223, 221, 221, 225, 135, 217, 226, 226, 226, 224, 226, 226, 228, 228, 226, 227, 227, 229, 230, 227, 229, 230, 229, 230, 230, 228, 229, 229, 231, 230, 229, 229, 229, 230, 230, 231, 229, 229, 229, 231, 231, 229, 229, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 230, 230, 231, 230, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 230, 231, 230, 230, 231, 232, 232, 231, 230, 231, 232, 232, 231, 230, 229, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 232, 233, 233, 232, 232, 232, 233, 234, 234, 234, 233, 233, 232, 209, 186, 185, 188, 189, 186, 188, 188, 183, 180, 184, 184, 189, 182, 186, 186, 193, 186, 194, 198, 204, 213, 223, 212, 191, 224, 191, 69, 43, 38, 41, 41, 46, 55, 67, 58, 47, 44, 40, 46, 40, 39, 43, 40, 40, 40, 41, 40, 43, 45, 50, 79, 49, 96, 64, 114, 160, 142, 54, 53, 48, 51, 50, 51, 51, 53, 52, 49, 54, 55, 76, 88, 66, 52, 56, 57, 71, 85, 130, 227, 234, 233, 229, 214, 163, 102, 71, 72, 88, 118, 167, 222, 230, 231, 229, 230, 229, 230, 231, 230, 231, 230, 230, 230, 232, 231, 231, 229, 230, 230, 231, 231, 229, 228, 229, 230, 230, 229, 226, 228, 224, 222, 224, 222, 219, 224, 132, 219, 227, 227, 227, 225, 225, 226, 228, 228, 226, 226, 228, 228, 229, 228, 228, 228, 229, 230, 230, 229, 228, 229, 230, 229, 229, 228, 230, 230, 230, 230, 229, 229, 229, 231, 230, 229, 229, 228, 230, 230, 231, 230, 229, 230, 231, 231, 230, 229, 230, 230, 231, 230, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 232, 231, 230, 230, 232, 231, 231, 231, 230, 230, 232, 231, 230, 230, 230, 231, 231, 232, 231, 230, 231, 231, 231, 231, 231, 230, 231, 231, 231, 231, 230, 231, 232, 231, 231, 231, 231, 232, 232, 232, 231, 232, 232, 233, 233, 232, 232, 232, 234, 233, 234, 234, 233, 233, 232, 218, 188, 184, 188, 190, 184, 189, 188, 181, 177, 178, 179, 183, 185, 188, 186, 188, 183, 188, 191, 201, 212, 224, 222, 193, 217, 205, 102, 39, 36, 39, 47, 100, 130, 94, 88, 101, 69, 40, 41, 39, 39, 39, 44, 41, 43, 44, 37, 40, 52, 47, 49, 50, 68, 60, 61, 144, 156, 80, 49, 47, 54, 47, 51, 50, 45, 49, 53, 55, 77, 131, 159, 103, 55, 52, 67, 73, 88, 139, 229, 234, 233, 227, 206, 148, 93, 67, 75, 98, 131, 172, 224, 230, 231, 230, 230, 229, 228, 230, 230, 231, 230, 230, 230, 231, 231, 231, 229, 231, 230, 230, 230, 229, 228, 228, 230, 230, 229, 228, 229, 227, 222, 226, 221, 217, 223, 123, 220, 228, 227, 227, 224, 227, 228, 228, 228, 226, 225, 225, 227, 228, 227, 228, 228, 229, 230, 229, 229, 228, 229, 229, 230, 228, 228, 229, 230, 231, 230, 229, 229, 229, 230, 231, 229, 229, 229, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 229, 229, 231, 232, 231, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 231, 230, 230, 231, 231, 232, 230, 230, 230, 232, 232, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 231, 230, 230, 231, 232, 232, 231, 231, 230, 232, 232, 232, 231, 231, 232, 233, 233, 232, 233, 232, 234, 234, 233, 233, 233, 233, 232, 221, 197, 181, 188, 190, 183, 191, 191, 181, 180, 176, 181, 184, 187, 188, 185, 186, 183, 186, 186, 199, 207, 221, 224, 202, 204, 220, 145, 41, 38, 48, 60, 153, 80, 48, 49, 73, 134, 45, 41, 37, 38, 39, 39, 42, 40, 44, 43, 40, 61, 53, 42, 46, 46, 57, 63, 96, 157, 129, 53, 46, 51, 47, 47, 48, 48, 51, 56, 56, 102, 119, 162, 99, 57, 52, 63, 69, 94, 157, 231, 233, 232, 228, 199, 145, 83, 70, 83, 107, 138, 181, 225, 230, 231, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 229, 230, 230, 229, 229, 228, 229, 230, 231, 230, 228, 228, 227, 222, 224, 221, 220, 223, 124, 220, 227, 226, 226, 226, 228, 228, 228, 227, 226, 226, 227, 228, 227, 227, 228, 229, 229, 229, 230, 229, 229, 230, 230, 232, 229, 227, 229, 230, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 231, 230, 230, 230, 230, 230, 232, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 232, 231, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 232, 230, 230, 229, 231, 231, 231, 230, 230, 230, 232, 232, 231, 231, 230, 232, 232, 232, 231, 232, 232, 233, 233, 232, 232, 233, 234, 234, 234, 233, 234, 233, 232, 223, 201, 185, 184, 190, 184, 190, 189, 186, 185, 177, 178, 184, 188, 189, 183, 184, 176, 173, 181, 196, 206, 216, 225, 211, 188, 223, 170, 63, 45, 52, 72, 161, 105, 47, 52, 61, 148, 46, 37, 37, 38, 36, 37, 43, 44, 40, 42, 36, 43, 40, 42, 41, 56, 74, 63, 61, 141, 155, 71, 48, 49, 56, 50, 46, 51, 50, 63, 75, 106, 105, 164, 114, 62, 54, 70, 74, 97, 176, 232, 233, 232, 227, 199, 150, 84, 76, 87, 118, 135, 187, 226, 230, 231, 231, 231, 230, 230, 230, 231, 231, 229, 230, 230, 230, 231, 231, 230, 230, 230, 230, 229, 229, 228, 230, 230, 231, 231, 229, 229, 227, 222, 226, 221, 221, 223, 126, 219, 225, 227, 224, 227, 225, 229, 227, 226, 228, 227, 228, 229, 228, 228, 229, 229, 229, 229, 230, 229, 230, 230, 230, 230, 229, 229, 230, 230, 230, 230, 229, 229, 230, 230, 231, 230, 230, 229, 231, 231, 231, 230, 230, 230, 231, 230, 230, 229, 229, 231, 231, 231, 229, 229, 230, 231, 231, 231, 229, 230, 231, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 230, 229, 231, 231, 231, 231, 230, 230, 230, 232, 231, 231, 230, 230, 232, 232, 231, 230, 229, 230, 232, 232, 230, 230, 229, 231, 232, 231, 230, 230, 231, 231, 232, 231, 231, 231, 232, 232, 232, 231, 231, 232, 233, 233, 232, 233, 232, 233, 234, 234, 233, 234, 233, 233, 227, 200, 187, 184, 189, 186, 188, 190, 186, 179, 177, 178, 176, 179, 179, 178, 172, 173, 168, 174, 189, 204, 216, 228, 217, 187, 207, 195, 101, 41, 46, 61, 162, 166, 120, 78, 111, 109, 39, 37, 42, 37, 32, 37, 34, 41, 41, 43, 49, 79, 84, 48, 44, 69, 87, 66, 72, 119, 161, 125, 67, 52, 48, 48, 48, 51, 56, 61, 117, 87, 88, 169, 127, 58, 57, 66, 76, 99, 196, 232, 232, 231, 226, 195, 151, 83, 78, 102, 119, 144, 198, 227, 230, 231, 231, 231, 230, 229, 231, 231, 232, 229, 230, 231, 231, 231, 230, 230, 230, 230, 230, 230, 229, 229, 229, 229, 230, 230, 229, 228, 227, 222, 226, 220, 221, 224, 125, 217, 225, 227, 225, 227, 226, 229, 227, 228, 227, 227, 229, 228, 228, 228, 228, 229, 229, 229, 229, 228, 228, 230, 231, 231, 230, 229, 229, 230, 229, 231, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 230, 230, 230, 229, 229, 230, 231, 231, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 232, 230, 230, 230, 231, 231, 231, 230, 229, 231, 231, 231, 230, 230, 230, 231, 232, 232, 231, 230, 231, 231, 232, 230, 229, 230, 231, 231, 231, 231, 230, 231, 232, 232, 231, 230, 231, 232, 232, 232, 231, 231, 232, 233, 233, 232, 233, 233, 233, 234, 235, 234, 234, 234, 232, 230, 198, 180, 180, 188, 188, 186, 192, 188, 181, 169, 172, 174, 169, 174, 172, 169, 170, 169, 173, 181, 200, 214, 224, 225, 195, 194, 205, 143, 47, 41, 50, 104, 171, 173, 164, 136, 67, 43, 39, 39, 36, 38, 46, 40, 40, 37, 39, 38, 51, 50, 40, 44, 53, 61, 52, 61, 73, 164, 163, 138, 55, 49, 42, 46, 52, 56, 75, 145, 83, 76, 161, 139, 59, 56, 64, 81, 101, 214, 233, 232, 230, 225, 185, 142, 77, 80, 113, 132, 149, 209, 228, 230, 231, 231, 230, 230, 229, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 229, 230, 229, 228, 228, 228, 230, 231, 231, 229, 229, 227, 222, 229, 221, 222, 224, 120, 216, 226, 227, 225, 227, 228, 229, 229, 227, 227, 227, 229, 227, 229, 229, 228, 228, 229, 229, 230, 228, 227, 230, 230, 230, 230, 228, 229, 231, 230, 230, 229, 229, 229, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 228, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 231, 230, 230, 230, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 232, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 232, 231, 231, 230, 232, 232, 232, 231, 232, 231, 232, 233, 232, 232, 232, 234, 234, 235, 234, 234, 234, 233, 231, 197, 185, 181, 189, 191, 188, 191, 190, 181, 171, 169, 164, 166, 166, 170, 171, 175, 170, 172, 177, 193, 209, 219, 222, 207, 183, 203, 177, 85, 44, 53, 136, 119, 124, 168, 172, 156, 92, 43, 34, 36, 33, 62, 43, 40, 42, 44, 42, 36, 43, 38, 41, 45, 40, 47, 56, 81, 164, 169, 133, 49, 45, 44, 51, 55, 61, 122, 159, 78, 72, 157, 143, 66, 80, 68, 92, 122, 225, 233, 231, 228, 221, 174, 129, 81, 97, 114, 133, 151, 211, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 231, 230, 231, 231, 231, 230, 229, 229, 230, 229, 228, 229, 227, 231, 231, 229, 229, 230, 228, 221, 226, 224, 223, 224, 127, 220, 225, 226, 225, 228, 227, 228, 229, 228, 226, 227, 228, 228, 229, 227, 228, 228, 229, 230, 229, 228, 228, 228, 230, 230, 229, 228, 229, 230, 230, 231, 229, 229, 229, 231, 231, 230, 230, 230, 231, 231, 231, 229, 229, 230, 231, 231, 230, 230, 229, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 232, 232, 231, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 231, 230, 231, 231, 232, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 230, 228, 230, 231, 231, 231, 231, 230, 230, 232, 232, 231, 231, 231, 232, 232, 232, 231, 232, 232, 232, 233, 233, 232, 232, 233, 234, 234, 234, 234, 234, 234, 232, 211, 188, 181, 186, 192, 190, 195, 191, 190, 181, 167, 162, 160, 170, 166, 168, 173, 170, 166, 177, 189, 206, 212, 221, 216, 193, 192, 200, 139, 54, 100, 151, 52, 54, 70, 118, 159, 151, 49, 38, 40, 39, 40, 38, 36, 39, 42, 45, 38, 74, 38, 46, 39, 42, 47, 53, 87, 124, 185, 181, 60, 53, 53, 55, 58, 67, 139, 143, 86, 76, 154, 154, 94, 85, 76, 92, 162, 229, 232, 231, 227, 213, 166, 119, 85, 105, 120, 136, 156, 218, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 231, 229, 231, 231, 230, 230, 229, 229, 230, 229, 227, 229, 228, 231, 231, 230, 230, 230, 227, 222, 229, 226, 221, 223, 121, 216, 225, 226, 226, 227, 228, 229, 229, 228, 228, 227, 229, 229, 227, 228, 228, 228, 229, 230, 229, 228, 229, 228, 230, 230, 229, 229, 229, 230, 231, 231, 229, 230, 230, 231, 231, 230, 230, 229, 230, 230, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 231, 229, 229, 230, 231, 231, 231, 230, 230, 230, 231, 232, 231, 231, 231, 232, 232, 232, 232, 231, 232, 233, 233, 232, 232, 232, 233, 234, 234, 234, 234, 234, 234, 232, 222, 196, 183, 186, 188, 189, 193, 193, 194, 183, 169, 162, 163, 168, 171, 167, 169, 166, 172, 175, 179, 199, 211, 215, 219, 206, 185, 212, 178, 90, 115, 148, 43, 43, 41, 53, 104, 162, 66, 41, 42, 45, 46, 46, 46, 42, 41, 39, 38, 41, 47, 48, 44, 60, 40, 57, 52, 59, 163, 205, 113, 71, 68, 76, 79, 82, 81, 63, 58, 56, 148, 156, 68, 65, 78, 105, 190, 232, 231, 230, 226, 195, 159, 98, 103, 115, 124, 138, 176, 221, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 230, 231, 231, 229, 229, 229, 230, 230, 229, 228, 229, 230, 231, 229, 229, 230, 227, 222, 228, 222, 218, 224, 117, 220, 226, 226, 227, 225, 227, 229, 228, 227, 227, 226, 228, 228, 228, 227, 227, 228, 229, 230, 229, 229, 228, 229, 230, 230, 229, 229, 229, 230, 230, 230, 230, 229, 230, 231, 231, 229, 229, 230, 231, 230, 230, 229, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 229, 229, 230, 231, 232, 231, 230, 230, 231, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 230, 230, 230, 231, 231, 230, 229, 230, 230, 231, 232, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 232, 231, 231, 230, 232, 232, 232, 231, 231, 232, 233, 233, 233, 232, 232, 233, 234, 234, 233, 234, 234, 234, 232, 227, 206, 185, 180, 190, 192, 194, 197, 196, 185, 171, 164, 161, 164, 175, 168, 172, 162, 164, 169, 172, 189, 202, 208, 218, 213, 193, 197, 195, 144, 95, 149, 56, 34, 38, 48, 70, 155, 58, 80, 137, 142, 149, 142, 138, 135, 104, 35, 35, 39, 52, 61, 34, 66, 42, 67, 43, 61, 96, 204, 173, 149, 167, 163, 168, 160, 143, 56, 53, 55, 140, 164, 69, 64, 110, 184, 223, 232, 231, 227, 224, 182, 147, 94, 110, 123, 134, 146, 190, 224, 230, 230, 231, 230, 230, 230, 229, 231, 231, 231, 230, 230, 230, 231, 231, 231, 229, 229, 229, 230, 231, 228, 228, 229, 230, 231, 230, 230, 230, 227, 222, 228, 222, 222, 224, 119, 217, 225, 226, 227, 226, 227, 228, 228, 227, 228, 227, 228, 229, 230, 228, 227, 227, 229, 229, 230, 228, 228, 229, 230, 231, 229, 229, 229, 230, 231, 231, 230, 230, 229, 231, 230, 230, 229, 230, 231, 230, 230, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 229, 229, 230, 231, 232, 230, 230, 230, 231, 232, 231, 230, 230, 230, 232, 231, 231, 230, 230, 231, 231, 231, 231, 230, 230, 231, 231, 231, 229, 230, 230, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 230, 232, 232, 232, 231, 231, 232, 233, 232, 232, 232, 232, 233, 234, 234, 233, 234, 234, 235, 233, 230, 211, 185, 177, 188, 193, 192, 195, 200, 191, 177, 164, 162, 170, 174, 177, 169, 169, 157, 145, 173, 177, 191, 205, 221, 218, 202, 182, 196, 177, 98, 125, 114, 50, 38, 44, 103, 105, 46, 122, 173, 179, 182, 180, 174, 164, 92, 40, 42, 41, 42, 39, 43, 63, 51, 46, 39, 51, 62, 169, 201, 152, 156, 149, 150, 133, 105, 50, 51, 58, 120, 137, 66, 71, 95, 172, 229, 232, 231, 226, 214, 173, 131, 98, 116, 124, 135, 144, 205, 227, 230, 230, 231, 231, 230, 230, 230, 230, 231, 232, 230, 230, 230, 231, 231, 230, 228, 228, 228, 230, 231, 229, 229, 228, 230, 231, 231, 229, 229, 228, 223, 228, 224, 222, 226, 114, 217, 225, 226, 228, 226, 228, 226, 227, 227, 227, 228, 228, 229, 230, 228, 227, 227, 230, 230, 230, 228, 228, 229, 230, 229, 229, 228, 229, 231, 230, 231, 229, 230, 230, 231, 231, 230, 229, 229, 231, 231, 230, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 230, 231, 230, 230, 229, 229, 231, 231, 231, 230, 230, 232, 232, 231, 230, 230, 231, 231, 231, 231, 230, 230, 231, 231, 231, 231, 230, 231, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 231, 231, 229, 232, 232, 232, 231, 231, 231, 232, 232, 232, 232, 232, 232, 234, 234, 233, 233, 234, 234, 234, 230, 214, 185, 184, 188, 191, 191, 200, 205, 191, 182, 167, 166, 166, 177, 186, 175, 174, 173, 164, 176, 181, 186, 202, 213, 218, 210, 190, 187, 186, 145, 70, 94, 89, 70, 71, 72, 43, 43, 84, 93, 100, 100, 98, 98, 142, 48, 41, 41, 38, 46, 89, 119, 98, 127, 118, 59, 50, 59, 119, 198, 135, 70, 79, 73, 62, 53, 49, 43, 48, 52, 58, 63, 73, 94, 204, 231, 230, 228, 222, 198, 159, 114, 107, 120, 130, 136, 162, 216, 229, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 231, 230, 230, 231, 231, 230, 229, 229, 228, 230, 230, 228, 229, 229, 231, 231, 231, 230, 229, 227, 222, 226, 223, 222, 224, 116, 214, 225, 226, 226, 225, 224, 228, 228, 228, 226, 227, 228, 230, 230, 229, 228, 229, 229, 230, 230, 227, 228, 229, 230, 230, 229, 228, 230, 231, 230, 231, 229, 230, 229, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 229, 229, 230, 231, 231, 230, 229, 230, 231, 231, 230, 230, 230, 231, 230, 231, 230, 230, 230, 231, 231, 231, 231, 230, 230, 232, 232, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 231, 230, 230, 230, 230, 232, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 230, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 232, 232, 233, 234, 234, 233, 233, 233, 235, 233, 230, 222, 181, 182, 181, 192, 194, 194, 201, 194, 185, 171, 167, 167, 178, 187, 184, 181, 178, 181, 183, 189, 183, 193, 206, 215, 216, 208, 181, 196, 175, 114, 47, 41, 41, 36, 36, 38, 35, 38, 37, 38, 46, 53, 119, 112, 39, 37, 44, 48, 91, 140, 60, 52, 75, 145, 131, 51, 50, 64, 163, 149, 104, 95, 107, 127, 83, 54, 42, 49, 50, 54, 65, 83, 146, 222, 232, 230, 224, 217, 173, 141, 118, 116, 126, 128, 139, 182, 224, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 231, 230, 230, 230, 230, 230, 230, 230, 229, 229, 230, 230, 228, 229, 229, 231, 231, 230, 228, 229, 227, 223, 227, 225, 222, 224, 113, 210, 227, 226, 225, 222, 226, 228, 228, 226, 228, 227, 227, 229, 229, 228, 227, 228, 229, 229, 230, 228, 228, 229, 229, 230, 228, 228, 230, 231, 230, 230, 230, 229, 230, 231, 230, 229, 230, 229, 231, 231, 230, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 231, 230, 230, 230, 231, 232, 231, 229, 230, 230, 231, 232, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 232, 231, 231, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 233, 233, 233, 233, 233, 233, 234, 234, 232, 228, 186, 181, 185, 186, 195, 192, 197, 199, 192, 176, 166, 162, 177, 188, 185, 184, 185, 186, 183, 191, 187, 188, 199, 211, 212, 215, 189, 185, 194, 159, 79, 42, 37, 37, 33, 36, 34, 38, 38, 43, 52, 81, 156, 74, 35, 36, 53, 58, 147, 121, 43, 48, 47, 106, 114, 48, 46, 47, 58, 95, 50, 51, 58, 108, 151, 84, 45, 51, 48, 58, 75, 88, 197, 228, 230, 228, 224, 194, 157, 127, 117, 117, 122, 129, 147, 201, 228, 229, 230, 230, 231, 232, 231, 230, 230, 231, 232, 231, 229, 230, 229, 230, 230, 230, 230, 230, 229, 229, 228, 229, 229, 229, 230, 230, 230, 230, 229, 227, 224, 225, 225, 223, 223, 114, 213, 226, 227, 224, 224, 225, 227, 227, 226, 227, 228, 228, 229, 228, 227, 228, 228, 230, 230, 230, 229, 230, 229, 229, 230, 230, 229, 229, 230, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 230, 231, 231, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 229, 231, 231, 231, 230, 230, 230, 231, 231, 231, 229, 230, 231, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 232, 230, 230, 231, 232, 233, 231, 231, 231, 232, 233, 233, 233, 232, 234, 234, 234, 232, 227, 204, 178, 183, 189, 193, 190, 192, 196, 193, 183, 170, 170, 178, 186, 183, 183, 184, 190, 185, 184, 190, 180, 189, 206, 204, 205, 206, 184, 188, 184, 146, 63, 38, 37, 32, 35, 38, 35, 35, 40, 55, 134, 156, 48, 37, 40, 50, 89, 168, 93, 40, 41, 45, 52, 48, 41, 42, 40, 53, 97, 43, 45, 56, 67, 155, 137, 51, 48, 56, 60, 82, 140, 223, 227, 228, 225, 217, 170, 142, 121, 121, 118, 124, 137, 168, 217, 230, 230, 229, 230, 232, 231, 231, 230, 230, 230, 231, 231, 229, 229, 230, 231, 230, 230, 229, 229, 227, 229, 229, 228, 227, 228, 230, 229, 230, 228, 229, 226, 222, 229, 225, 222, 224, 121, 214, 226, 227, 227, 226, 227, 228, 227, 228, 228, 227, 228, 230, 228, 227, 228, 227, 230, 229, 230, 230, 229, 228, 229, 230, 230, 229, 229, 230, 230, 231, 230, 229, 230, 231, 231, 230, 230, 229, 230, 231, 231, 230, 229, 230, 231, 231, 231, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 229, 230, 231, 230, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 232, 231, 230, 230, 229, 231, 231, 230, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 232, 231, 231, 230, 231, 231, 232, 231, 231, 230, 231, 232, 233, 232, 232, 231, 233, 234, 233, 233, 233, 233, 235, 235, 233, 228, 223, 177, 185, 183, 194, 191, 193, 199, 193, 189, 176, 168, 174, 181, 182, 186, 189, 190, 192, 191, 189, 189, 182, 191, 202, 206, 211, 197, 176, 192, 176, 131, 50, 39, 35, 36, 35, 36, 39, 51, 68, 165, 137, 37, 35, 39, 47, 123, 166, 77, 42, 61, 84, 98, 63, 41, 41, 47, 104, 115, 40, 42, 51, 57, 145, 158, 67, 52, 62, 71, 101, 203, 227, 226, 227, 224, 192, 161, 127, 122, 118, 118, 123, 137, 191, 226, 231, 229, 229, 229, 230, 231, 230, 230, 230, 230, 232, 230, 230, 229, 228, 230, 230, 230, 229, 228, 227, 229, 228, 228, 228, 227, 228, 229, 229, 229, 229, 225, 221, 227, 224, 223, 225, 131, 213, 225, 229, 225, 225, 226, 227, 228, 228, 228, 227, 227, 229, 228, 227, 226, 225, 225, 228, 228, 228, 229, 228, 229, 229, 229, 229, 228, 230, 230, 230, 230, 229, 230, 231, 231, 230, 228, 229, 230, 231, 231, 229, 229, 229, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 229, 229, 230, 231, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 229, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 231, 232, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 232, 231, 233, 233, 233, 232, 232, 233, 234, 235, 233, 231, 228, 191, 180, 186, 184, 192, 192, 192, 192, 193, 179, 173, 175, 182, 184, 184, 189, 186, 189, 186, 189, 188, 184, 182, 196, 208, 211, 208, 191, 178, 189, 172, 114, 47, 37, 37, 34, 41, 35, 47, 108, 165, 109, 37, 34, 38, 46, 132, 165, 72, 54, 67, 73, 121, 142, 102, 43, 45, 115, 84, 40, 41, 49, 55, 143, 160, 69, 54, 64, 86, 173, 221, 226, 225, 225, 210, 175, 133, 121, 119, 115, 117, 123, 158, 209, 229, 230, 230, 229, 228, 230, 231, 230, 229, 230, 229, 232, 231, 229, 229, 227, 229, 230, 230, 229, 228, 228, 228, 229, 227, 225, 225, 228, 228, 227, 229, 228, 224, 220, 227, 224, 224, 224, 126, 214, 226, 228, 225, 227, 227, 227, 229, 229, 228, 227, 227, 229, 228, 226, 223, 224, 227, 228, 228, 228, 227, 227, 227, 228, 228, 227, 229, 230, 230, 229, 230, 229, 230, 230, 230, 230, 230, 230, 230, 231, 231, 229, 229, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 231, 232, 231, 231, 230, 230, 230, 231, 231, 230, 231, 231, 231, 231, 231, 231, 231, 231, 232, 232, 231, 231, 231, 232, 233, 232, 231, 231, 232, 233, 233, 233, 233, 232, 234, 234, 234, 232, 228, 217, 177, 185, 182, 191, 191, 192, 198, 192, 188, 175, 173, 179, 182, 184, 186, 188, 184, 187, 187, 184, 186, 178, 186, 202, 205, 209, 203, 183, 179, 193, 163, 109, 42, 35, 35, 39, 41, 43, 141, 169, 96, 34, 37, 40, 49, 136, 166, 84, 56, 42, 44, 53, 135, 158, 77, 50, 92, 94, 41, 41, 50, 54, 142, 160, 69, 62, 76, 138, 216, 227, 225, 224, 218, 177, 158, 121, 111, 112, 106, 107, 126, 180, 220, 230, 231, 229, 228, 229, 230, 231, 230, 229, 229, 229, 230, 231, 228, 229, 227, 228, 229, 228, 228, 226, 225, 228, 228, 226, 224, 225, 227, 229, 229, 228, 227, 224, 219, 225, 225, 224, 225, 135, 220, 227, 225, 225, 227, 228, 228, 229, 230, 229, 227, 226, 228, 227, 224, 223, 224, 224, 228, 229, 227, 224, 226, 225, 224, 225, 227, 228, 230, 230, 228, 229, 229, 230, 230, 230, 230, 230, 230, 231, 231, 231, 229, 229, 229, 231, 231, 231, 229, 230, 231, 232, 231, 230, 230, 230, 231, 231, 231, 229, 230, 230, 230, 231, 230, 230, 230, 230, 231, 232, 230, 230, 230, 231, 230, 229, 229, 230, 230, 230, 230, 230, 230, 230, 232, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 231, 230, 230, 232, 232, 231, 230, 230, 232, 232, 231, 230, 231, 231, 232, 232, 232, 231, 231, 233, 233, 233, 233, 232, 233, 234, 234, 234, 231, 230, 227, 187, 183, 183, 187, 187, 195, 189, 192, 190, 182, 171, 178, 178, 180, 187, 187, 185, 187, 192, 185, 185, 181, 173, 193, 204, 209, 208, 201, 179, 184, 189, 162, 100, 42, 36, 36, 44, 46, 154, 167, 73, 37, 33, 41, 48, 132, 169, 87, 59, 36, 41, 46, 94, 161, 123, 45, 50, 98, 41, 41, 56, 71, 154, 129, 58, 73, 119, 208, 224, 226, 224, 220, 191, 165, 125, 111, 97, 103, 100, 109, 144, 211, 228, 231, 230, 229, 228, 229, 229, 229, 230, 228, 229, 228, 231, 229, 228, 227, 226, 229, 229, 227, 225, 224, 226, 226, 226, 225, 225, 226, 226, 226, 227, 226, 226, 222, 218, 227, 224, 222, 226, 127, 218, 228, 226, 225, 226, 227, 229, 229, 230, 228, 228, 227, 228, 225, 223, 221, 222, 223, 227, 227, 225, 224, 226, 226, 225, 225, 227, 226, 228, 227, 227, 227, 227, 229, 230, 231, 230, 229, 230, 231, 231, 231, 229, 229, 229, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 230, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 230, 229, 230, 230, 230, 231, 229, 229, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 231, 229, 230, 231, 231, 231, 230, 230, 230, 231, 232, 231, 231, 230, 231, 231, 231, 231, 231, 231, 232, 232, 232, 231, 232, 233, 233, 233, 232, 232, 233, 234, 234, 233, 232, 231, 228, 212, 183, 184, 181, 186, 194, 191, 193, 194, 188, 174, 179, 180, 182, 184, 187, 186, 188, 186, 185, 178, 180, 168, 179, 194, 197, 207, 209, 199, 178, 174, 185, 159, 101, 47, 41, 48, 53, 159, 163, 68, 34, 37, 36, 50, 112, 160, 104, 60, 36, 37, 51, 72, 156, 144, 45, 41, 68, 90, 69, 70, 128, 135, 67, 71, 112, 196, 220, 223, 224, 219, 197, 164, 129, 116, 88, 87, 87, 89, 110, 179, 220, 229, 230, 230, 229, 228, 229, 229, 229, 230, 228, 228, 229, 230, 230, 227, 228, 228, 230, 225, 225, 222, 225, 227, 226, 227, 226, 224, 224, 227, 225, 225, 223, 222, 220, 215, 228, 224, 223, 223, 119, 217, 227, 227, 225, 227, 227, 229, 228, 229, 228, 226, 226, 227, 225, 220, 221, 224, 225, 225, 229, 226, 225, 226, 224, 226, 225, 225, 225, 227, 227, 228, 227, 229, 228, 228, 230, 230, 228, 228, 230, 230, 230, 229, 230, 230, 230, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 229, 230, 230, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 229, 230, 231, 230, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 232, 231, 230, 229, 231, 231, 232, 231, 230, 231, 232, 233, 231, 231, 231, 232, 233, 233, 232, 232, 233, 233, 233, 233, 232, 232, 230, 227, 180, 182, 177, 184, 194, 189, 197, 191, 189, 182, 176, 174, 178, 181, 183, 188, 186, 184, 181, 172, 165, 156, 163, 174, 192, 202, 203, 205, 193, 173, 182, 178, 163, 111, 54, 53, 58, 151, 150, 60, 34, 36, 37, 52, 86, 157, 118, 74, 40, 40, 48, 60, 160, 149, 42, 38, 40, 50, 72, 77, 82, 84, 151, 117, 194, 218, 218, 220, 216, 196, 171, 128, 112, 90, 79, 76, 82, 91, 145, 206, 225, 230, 230, 230, 229, 228, 229, 230, 229, 229, 227, 229, 230, 230, 230, 226, 228, 227, 229, 225, 227, 226, 226, 225, 225, 226, 226, 223, 223, 226, 223, 225, 224, 222, 220, 214, 226, 224, 221, 225, 118, 220, 227, 227, 226, 229, 227, 227, 229, 228, 228, 226, 227, 224, 222, 217, 218, 220, 224, 225, 228, 225, 226, 224, 225, 224, 224, 226, 227, 226, 227, 228, 226, 229, 227, 228, 229, 229, 228, 229, 230, 228, 229, 229, 229, 229, 230, 230, 231, 229, 229, 230, 230, 231, 230, 230, 229, 231, 231, 229, 229, 229, 230, 230, 231, 229, 229, 230, 231, 231, 230, 230, 229, 230, 230, 230, 229, 229, 229, 230, 229, 229, 228, 228, 229, 230, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 232, 231, 230, 230, 231, 231, 231, 231, 230, 231, 232, 232, 232, 231, 231, 233, 233, 232, 232, 232, 232, 232, 233, 233, 233, 233, 232, 230, 205, 177, 182, 178, 191, 195, 193, 187, 190, 188, 181, 168, 175, 178, 179, 187, 187, 185, 176, 162, 154, 151, 154, 162, 178, 190, 202, 208, 203, 192, 171, 175, 183, 166, 134, 111, 82, 57, 53, 40, 32, 34, 36, 51, 53, 142, 142, 74, 56, 44, 49, 57, 155, 129, 37, 40, 39, 36, 43, 46, 58, 102, 188, 200, 213, 219, 215, 216, 194, 173, 142, 104, 99, 69, 73, 74, 80, 117, 188, 221, 228, 230, 230, 230, 229, 229, 229, 230, 228, 229, 228, 229, 229, 230, 229, 227, 227, 226, 228, 224, 227, 225, 227, 226, 227, 227, 226, 222, 222, 225, 224, 226, 224, 223, 221, 214, 226, 224, 221, 224, 121, 219, 225, 225, 227, 227, 227, 229, 230, 226, 226, 224, 226, 224, 226, 218, 217, 220, 224, 224, 225, 224, 224, 225, 226, 225, 223, 227, 225, 227, 228, 227, 227, 227, 227, 228, 229, 229, 229, 229, 230, 229, 230, 228, 229, 229, 229, 231, 230, 229, 229, 230, 230, 229, 229, 229, 228, 229, 228, 227, 226, 227, 227, 227, 227, 224, 226, 224, 224, 223, 220, 218, 217, 214, 217, 210, 206, 208, 203, 198, 199, 196, 189, 189, 190, 199, 219, 221, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 231, 230, 231, 231, 231, 231, 230, 230, 231, 231, 231, 231, 231, 231, 232, 232, 231, 231, 231, 232, 233, 233, 232, 232, 232, 233, 234, 234, 233, 233, 232, 230, 227, 171, 176, 179, 184, 193, 193, 186, 188, 186, 185, 175, 167, 174, 178, 185, 184, 179, 176, 153, 149, 149, 146, 146, 160, 175, 192, 199, 204, 199, 192, 168, 176, 183, 177, 153, 103, 50, 43, 41, 35, 36, 38, 44, 52, 99, 137, 85, 57, 41, 52, 72, 153, 77, 34, 38, 35, 36, 44, 54, 78, 157, 205, 215, 215, 210, 205, 189, 164, 129, 105, 91, 74, 68, 65, 74, 96, 166, 215, 227, 229, 231, 230, 230, 228, 228, 229, 229, 229, 229, 228, 229, 229, 230, 227, 228, 227, 226, 226, 227, 227, 224, 227, 228, 229, 228, 226, 225, 224, 224, 225, 224, 225, 223, 220, 212, 229, 226, 223, 227, 131, 223, 225, 228, 227, 228, 229, 231, 231, 228, 223, 210, 203, 198, 202, 193, 194, 193, 195, 196, 196, 194, 196, 193, 196, 197, 197, 200, 197, 200, 204, 199, 202, 206, 204, 206, 206, 208, 210, 211, 211, 212, 219, 214, 215, 218, 218, 226, 212, 203, 201, 198, 193, 189, 186, 182, 178, 169, 166, 159, 160, 163, 157, 152, 156, 148, 148, 136, 138, 134, 133, 133, 128, 122, 126, 116, 117, 116, 111, 111, 115, 120, 124, 124, 132, 154, 132, 140, 226, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 231, 231, 230, 230, 231, 232, 231, 231, 231, 231, 232, 232, 231, 231, 231, 232, 233, 232, 231, 232, 232, 233, 234, 234, 233, 234, 234, 233, 228, 201, 172, 178, 182, 190, 189, 185, 185, 188, 184, 181, 173, 164, 175, 182, 183, 184, 171, 153, 146, 142, 135, 139, 140, 150, 171, 189, 193, 199, 203, 190, 172, 172, 186, 186, 167, 123, 68, 50, 42, 39, 44, 39, 46, 66, 98, 131, 62, 48, 51, 109, 118, 39, 37, 36, 39, 43, 59, 111, 175, 202, 208, 209, 206, 199, 178, 161, 130, 105, 100, 66, 69, 71, 62, 85, 143, 203, 226, 228, 229, 230, 231, 229, 229, 229, 230, 230, 230, 228, 229, 228, 227, 228, 228, 228, 227, 227, 227, 225, 223, 224, 226, 226, 227, 228, 224, 226, 225, 225, 224, 225, 225, 221, 218, 214, 233, 229, 226, 231, 134, 226, 234, 235, 235, 237, 237, 240, 238, 227, 204, 95, 91, 82, 80, 81, 81, 80, 85, 85, 85, 79, 82, 80, 81, 78, 82, 79, 77, 81, 83, 84, 81, 81, 82, 87, 86, 81, 88, 87, 92, 94, 103, 97, 101, 108, 127, 160, 143, 124, 131, 133, 124, 110, 109, 104, 97, 96, 99, 96, 95, 95, 92, 95, 99, 97, 93, 88, 95, 96, 93, 91, 90, 94, 89, 91, 91, 94, 97, 103, 107, 111, 112, 114, 110, 151, 106, 117, 225, 230, 231, 230, 231, 229, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 230, 232, 232, 230, 230, 231, 232, 232, 232, 231, 231, 232, 233, 232, 232, 232, 232, 234, 234, 233, 233, 233, 235, 233, 230, 224, 171, 178, 183, 182, 187, 191, 186, 188, 189, 187, 180, 168, 162, 167, 173, 173, 161, 139, 140, 131, 127, 131, 127, 138, 143, 171, 182, 188, 200, 199, 195, 177, 161, 176, 187, 177, 159, 108, 58, 45, 38, 48, 46, 52, 55, 95, 111, 96, 82, 93, 54, 55, 77, 90, 65, 97, 154, 187, 201, 201, 201, 201, 182, 170, 155, 125, 107, 100, 64, 59, 67, 69, 76, 131, 193, 221, 229, 229, 230, 231, 231, 230, 230, 229, 229, 230, 231, 230, 230, 228, 228, 230, 228, 225, 228, 227, 226, 225, 225, 223, 225, 227, 228, 225, 225, 226, 225, 224, 226, 223, 223, 223, 218, 215, 235, 229, 228, 232, 123, 226, 233, 232, 235, 236, 238, 240, 238, 228, 203, 84, 80, 70, 75, 72, 71, 69, 73, 76, 75, 71, 74, 72, 74, 72, 66, 67, 70, 69, 72, 75, 71, 76, 73, 75, 74, 73, 74, 70, 76, 78, 79, 75, 80, 99, 139, 158, 159, 130, 143, 121, 109, 95, 87, 92, 86, 86, 89, 88, 95, 86, 86, 90, 92, 89, 90, 86, 88, 91, 90, 79, 83, 80, 87, 86, 90, 95, 104, 112, 116, 124, 120, 146, 106, 145, 105, 118, 224, 230, 231, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 232, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 232, 232, 232, 233, 234, 233, 233, 233, 235, 235, 234, 229, 204, 177, 178, 187, 187, 190, 189, 187, 188, 188, 190, 178, 170, 155, 153, 148, 142, 143, 137, 132, 140, 123, 122, 121, 128, 138, 162, 174, 184, 191, 200, 195, 183, 163, 162, 178, 182, 171, 150, 110, 79, 95, 93, 88, 88, 84, 71, 170, 97, 109, 113, 131, 132, 138, 151, 175, 188, 190, 197, 191, 182, 174, 167, 146, 108, 120, 97, 64, 53, 61, 62, 75, 121, 185, 222, 230, 230, 229, 230, 231, 231, 230, 229, 229, 230, 231, 230, 229, 229, 228, 230, 229, 230, 226, 227, 228, 224, 225, 224, 224, 224, 228, 226, 226, 226, 225, 226, 226, 224, 222, 223, 221, 219, 213, 234, 229, 230, 230, 127, 224, 230, 233, 234, 235, 237, 241, 238, 228, 202, 87, 79, 98, 74, 69, 70, 73, 72, 73, 77, 74, 74, 75, 74, 73, 70, 68, 72, 70, 71, 75, 73, 74, 80, 80, 83, 80, 83, 80, 84, 84, 82, 79, 84, 96, 148, 170, 179, 166, 207, 113, 115, 103, 89, 97, 113, 103, 102, 133, 160, 165, 165, 171, 174, 173, 154, 150, 153, 167, 131, 102, 140, 129, 131, 143, 153, 160, 169, 170, 178, 176, 160, 158, 105, 139, 101, 116, 222, 230, 231, 231, 230, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 231, 231, 231, 230, 232, 232, 231, 230, 230, 230, 232, 232, 232, 231, 231, 232, 232, 232, 231, 232, 232, 234, 234, 233, 233, 233, 235, 235, 234, 231, 227, 191, 174, 181, 183, 184, 191, 192, 187, 189, 189, 183, 173, 157, 147, 142, 136, 135, 135, 133, 132, 129, 123, 114, 113, 118, 134, 158, 167, 181, 192, 195, 199, 189, 169, 157, 160, 178, 180, 164, 159, 139, 119, 110, 105, 107, 108, 150, 117, 128, 139, 153, 161, 165, 169, 172, 174, 176, 175, 171, 165, 151, 126, 119, 118, 90, 62, 53, 56, 59, 73, 117, 180, 217, 229, 231, 230, 230, 229, 231, 230, 231, 229, 229, 230, 231, 230, 229, 229, 227, 227, 228, 228, 226, 227, 228, 226, 227, 226, 225, 224, 225, 224, 224, 225, 224, 223, 224, 225, 224, 223, 222, 219, 218, 231, 228, 227, 228, 120, 221, 229, 231, 231, 233, 235, 236, 232, 223, 190, 89, 78, 151, 75, 75, 82, 121, 130, 138, 144, 153, 156, 168, 164, 159, 142, 141, 148, 156, 146, 152, 153, 141, 186, 191, 192, 193, 195, 194, 197, 192, 181, 158, 95, 92, 136, 170, 190, 169, 212, 190, 211, 183, 153, 147, 177, 158, 146, 200, 223, 225, 225, 225, 222, 217, 184, 192, 171, 162, 127, 108, 150, 144, 148, 160, 170, 168, 177, 176, 183, 180, 163, 155, 104, 143, 102, 112, 223, 229, 232, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 228, 230, 231, 232, 231, 230, 230, 231, 232, 232, 232, 231, 231, 232, 233, 232, 232, 232, 232, 234, 234, 233, 233, 233, 234, 235, 235, 233, 230, 225, 177, 177, 179, 180, 187, 192, 190, 187, 192, 187, 185, 174, 159, 144, 137, 133, 135, 128, 129, 133, 120, 117, 89, 81, 110, 154, 147, 156, 175, 188, 198, 193, 190, 185, 166, 153, 154, 167, 172, 170, 168, 161, 154, 147, 142, 153, 147, 142, 152, 156, 156, 160, 165, 169, 174, 172, 170, 155, 129, 125, 131, 116, 80, 63, 69, 61, 56, 68, 124, 182, 217, 227, 230, 231, 230, 229, 229, 229, 229, 229, 229, 230, 229, 230, 229, 230, 228, 228, 227, 229, 228, 226, 228, 227, 225, 227, 226, 224, 227, 226, 226, 225, 227, 226, 225, 226, 223, 224, 224, 223, 221, 219, 231, 227, 227, 228, 122, 221, 231, 231, 230, 233, 233, 236, 232, 223, 190, 87, 88, 105, 85, 96, 103, 177, 181, 182, 186, 185, 185, 187, 185, 159, 137, 141, 139, 143, 142, 144, 158, 176, 219, 222, 223, 223, 220, 222, 223, 214, 201, 187, 107, 94, 150, 176, 178, 164, 201, 200, 222, 195, 182, 172, 192, 171, 160, 208, 229, 231, 231, 232, 227, 217, 172, 151, 100, 85, 78, 79, 95, 126, 146, 155, 168, 171, 177, 180, 183, 179, 156, 158, 104, 136, 97, 121, 225, 230, 231, 231, 231, 230, 230, 229, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 230, 230, 230, 231, 232, 232, 231, 230, 231, 232, 232, 231, 231, 231, 231, 231, 232, 232, 232, 232, 233, 233, 233, 232, 233, 234, 235, 235, 234, 233, 230, 223, 200, 183, 183, 181, 188, 194, 190, 188, 187, 184, 180, 170, 160, 151, 135, 132, 132, 126, 130, 125, 126, 113, 79, 161, 155, 109, 119, 144, 168, 181, 186, 189, 192, 194, 184, 165, 145, 140, 152, 166, 171, 169, 178, 169, 168, 168, 172, 172, 173, 176, 173, 172, 166, 161, 146, 131, 136, 135, 135, 109, 69, 83, 60, 54, 64, 77, 119, 184, 219, 227, 230, 230, 230, 229, 228, 228, 229, 231, 230, 229, 229, 229, 229, 230, 229, 229, 229, 230, 228, 228, 227, 226, 223, 224, 227, 228, 225, 226, 228, 225, 226, 225, 225, 225, 225, 223, 223, 220, 223, 220, 216, 232, 228, 227, 228, 132, 224, 230, 232, 231, 234, 235, 237, 233, 222, 187, 87, 74, 94, 112, 119, 121, 130, 129, 131, 136, 134, 135, 140, 143, 146, 148, 152, 152, 141, 115, 125, 140, 174, 220, 226, 224, 224, 222, 222, 223, 220, 204, 192, 110, 87, 124, 176, 157, 160, 183, 203, 223, 203, 185, 183, 195, 179, 173, 207, 231, 232, 233, 233, 227, 213, 143, 80, 78, 85, 85, 79, 85, 102, 145, 158, 166, 172, 174, 180, 181, 182, 156, 159, 116, 142, 102, 122, 226, 230, 231, 231, 231, 229, 230, 230, 231, 231, 230, 230, 229, 231, 231, 231, 230, 230, 231, 231, 232, 230, 230, 230, 232, 232, 232, 231, 230, 231, 232, 232, 231, 231, 231, 231, 232, 233, 231, 232, 232, 233, 233, 232, 232, 232, 234, 235, 235, 234, 234, 233, 232, 226, 189, 182, 184, 183, 192, 195, 188, 182, 188, 185, 179, 171, 157, 145, 137, 131, 131, 127, 121, 124, 119, 77, 167, 116, 71, 79, 110, 126, 153, 168, 178, 186, 189, 190, 188, 180, 174, 164, 152, 143, 135, 142, 151, 159, 159, 158, 156, 162, 155, 148, 139, 135, 142, 149, 147, 145, 118, 79, 54, 45, 64, 79, 57, 63, 81, 141, 212, 227, 230, 230, 231, 232, 230, 229, 229, 230, 231, 230, 230, 229, 230, 230, 229, 229, 229, 229, 230, 230, 228, 225, 225, 222, 226, 228, 228, 226, 227, 226, 226, 227, 226, 224, 224, 225, 224, 224, 223, 224, 220, 218, 232, 227, 228, 227, 133, 224, 232, 233, 232, 235, 236, 236, 233, 222, 178, 94, 74, 87, 117, 125, 122, 122, 126, 137, 134, 138, 139, 145, 150, 151, 148, 151, 133, 117, 107, 119, 132, 179, 221, 227, 225, 222, 224, 216, 220, 221, 194, 189, 104, 86, 116, 181, 145, 171, 186, 205, 228, 226, 213, 190, 201, 195, 183, 210, 232, 233, 235, 233, 228, 209, 119, 76, 77, 85, 81, 79, 82, 94, 119, 154, 172, 174, 172, 180, 185, 185, 161, 172, 114, 144, 101, 124, 226, 230, 231, 231, 230, 229, 229, 230, 231, 230, 230, 230, 230, 232, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 231, 231, 232, 231, 231, 231, 232, 232, 233, 231, 231, 231, 233, 233, 232, 232, 232, 234, 234, 235, 234, 234, 234, 235, 233, 226, 192, 180, 185, 185, 189, 193, 184, 182, 181, 187, 183, 172, 163, 149, 142, 139, 126, 124, 116, 99, 99, 105, 45, 56, 52, 86, 94, 100, 129, 147, 164, 175, 180, 180, 185, 188, 183, 189, 179, 176, 166, 162, 155, 151, 152, 151, 156, 161, 168, 161, 162, 161, 153, 130, 100, 71, 55, 42, 46, 69, 76, 75, 65, 70, 123, 202, 226, 229, 230, 231, 231, 229, 228, 229, 229, 231, 230, 230, 229, 229, 230, 230, 230, 229, 229, 229, 227, 225, 224, 223, 221, 225, 227, 227, 225, 226, 227, 226, 226, 226, 225, 224, 223, 224, 222, 222, 223, 219, 215, 231, 228, 227, 228, 116, 218, 232, 232, 233, 234, 236, 236, 234, 222, 178, 89, 78, 81, 116, 127, 128, 128, 140, 141, 135, 138, 138, 147, 150, 144, 123, 91, 78, 83, 87, 100, 130, 184, 223, 224, 224, 224, 220, 220, 222, 216, 208, 194, 99, 92, 124, 200, 147, 171, 181, 214, 230, 230, 227, 220, 211, 205, 195, 219, 232, 233, 235, 233, 224, 207, 115, 91, 92, 87, 81, 74, 79, 83, 99, 151, 166, 178, 179, 182, 189, 184, 158, 173, 123, 150, 107, 122, 225, 230, 231, 231, 230, 229, 229, 230, 230, 231, 230, 229, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 231, 231, 231, 231, 232, 232, 233, 232, 231, 231, 232, 233, 233, 232, 232, 233, 234, 234, 233, 234, 234, 235, 235, 233, 228, 203, 184, 191, 185, 182, 186, 182, 176, 182, 179, 181, 174, 164, 154, 140, 127, 120, 116, 96, 172, 71, 52, 94, 104, 102, 95, 88, 90, 98, 116, 135, 150, 163, 168, 175, 180, 177, 179, 181, 179, 181, 182, 183, 176, 181, 177, 173, 172, 154, 142, 121, 98, 75, 66, 60, 67, 66, 60, 163, 137, 104, 102, 70, 86, 154, 213, 227, 229, 230, 230, 228, 229, 230, 230, 230, 230, 229, 228, 229, 229, 229, 228, 227, 228, 229, 229, 227, 225, 220, 219, 224, 227, 226, 225, 226, 226, 226, 227, 224, 224, 222, 222, 224, 220, 224, 223, 216, 214, 230, 229, 226, 229, 129, 225, 233, 232, 234, 234, 236, 237, 234, 223, 176, 86, 81, 86, 120, 120, 118, 110, 134, 140, 139, 135, 139, 149, 152, 133, 77, 73, 73, 75, 75, 86, 118, 189, 222, 224, 225, 224, 222, 220, 220, 220, 211, 197, 106, 94, 132, 203, 143, 171, 180, 217, 230, 231, 228, 228, 226, 215, 205, 221, 231, 231, 235, 232, 224, 214, 144, 178, 165, 129, 82, 71, 84, 82, 95, 149, 163, 179, 185, 181, 187, 183, 157, 172, 126, 158, 113, 120, 226, 230, 231, 231, 230, 229, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 230, 231, 232, 232, 232, 231, 231, 232, 232, 232, 232, 232, 232, 233, 234, 233, 233, 233, 234, 235, 236, 235, 233, 230, 214, 189, 187, 176, 178, 182, 181, 176, 176, 185, 183, 177, 166, 155, 138, 125, 109, 140, 152, 64, 55, 87, 98, 94, 89, 84, 83, 76, 78, 77, 95, 112, 124, 139, 150, 159, 163, 162, 166, 166, 168, 170, 165, 161, 147, 140, 121, 101, 84, 74, 70, 67, 70, 74, 89, 115, 126, 139, 153, 102, 128, 110, 73, 96, 172, 216, 228, 230, 231, 229, 229, 230, 230, 230, 231, 229, 228, 229, 229, 230, 228, 228, 227, 227, 227, 226, 224, 222, 220, 223, 225, 227, 225, 224, 227, 224, 225, 226, 224, 225, 223, 225, 224, 224, 221, 217, 212, 231, 227, 229, 230, 134, 228, 234, 233, 234, 235, 236, 238, 235, 224, 181, 85, 79, 82, 111, 107, 78, 76, 100, 124, 131, 140, 140, 143, 144, 103, 69, 68, 74, 74, 75, 81, 101, 186, 217, 222, 220, 221, 218, 212, 218, 220, 207, 199, 109, 90, 136, 200, 158, 172, 185, 217, 230, 228, 228, 229, 228, 227, 219, 222, 229, 228, 232, 231, 227, 216, 175, 189, 192, 175, 107, 78, 85, 86, 105, 160, 155, 169, 180, 184, 184, 178, 156, 166, 125, 154, 107, 128, 226, 229, 231, 231, 230, 230, 230, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 230, 230, 230, 231, 231, 231, 231, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 232, 232, 233, 232, 232, 232, 234, 233, 234, 233, 234, 234, 235, 236, 235, 235, 235, 232, 222, 191, 177, 148, 168, 180, 185, 177, 180, 182, 185, 185, 178, 161, 143, 122, 192, 94, 55, 63, 87, 87, 84, 80, 78, 73, 66, 67, 63, 70, 61, 63, 76, 79, 90, 100, 107, 108, 110, 113, 107, 94, 89, 76, 63, 51, 66, 70, 74, 86, 106, 129, 153, 180, 202, 200, 173, 148, 135, 88, 131, 99, 75, 105, 184, 221, 229, 230, 229, 228, 229, 228, 230, 230, 228, 228, 228, 229, 229, 227, 229, 227, 227, 228, 227, 224, 222, 221, 223, 225, 226, 226, 226, 225, 221, 224, 224, 223, 224, 223, 224, 224, 219, 219, 218, 214, 233, 230, 230, 231, 144, 229, 234, 233, 235, 236, 237, 238, 235, 222, 175, 80, 85, 76, 96, 97, 81, 86, 80, 94, 117, 128, 138, 144, 136, 84, 74, 66, 70, 70, 70, 77, 85, 173, 209, 210, 210, 209, 207, 200, 202, 199, 184, 180, 108, 87, 135, 204, 153, 168, 182, 208, 230, 228, 228, 229, 228, 229, 229, 228, 229, 231, 232, 231, 227, 211, 166, 152, 154, 175, 147, 88, 95, 96, 118, 161, 161, 167, 173, 172, 173, 160, 139, 171, 126, 152, 109, 130, 227, 229, 230, 230, 230, 230, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 231, 232, 233, 232, 232, 232, 234, 233, 234, 233, 232, 234, 235, 236, 235, 235, 236, 236, 234, 226, 198, 147, 126, 159, 181, 180, 179, 179, 178, 185, 180, 170, 132, 138, 162, 69, 59, 73, 99, 95, 90, 89, 93, 84, 75, 67, 69, 62, 54, 53, 55, 55, 52, 54, 55, 57, 57, 52, 56, 47, 44, 50, 56, 69, 74, 102, 155, 175, 191, 202, 213, 223, 227, 228, 216, 149, 150, 142, 94, 145, 85, 69, 118, 195, 224, 229, 229, 228, 229, 229, 230, 231, 228, 227, 228, 229, 229, 228, 227, 226, 227, 227, 226, 225, 222, 222, 223, 226, 226, 225, 227, 224, 223, 223, 224, 224, 223, 224, 222, 223, 221, 221, 219, 212, 232, 230, 228, 230, 130, 224, 233, 235, 235, 236, 236, 235, 234, 223, 169, 78, 78, 73, 79, 84, 124, 117, 99, 150, 192, 157, 160, 170, 155, 87, 92, 99, 103, 96, 88, 93, 98, 139, 164, 154, 145, 134, 125, 107, 98, 93, 79, 141, 104, 90, 134, 204, 157, 173, 182, 202, 229, 229, 230, 229, 230, 232, 231, 232, 231, 232, 232, 230, 226, 188, 126, 144, 126, 154, 176, 155, 127, 104, 146, 164, 160, 133, 133, 131, 136, 132, 122, 163, 126, 149, 109, 128, 226, 229, 231, 231, 230, 230, 230, 230, 231, 231, 230, 229, 230, 231, 232, 231, 230, 230, 229, 231, 231, 230, 230, 230, 231, 231, 230, 230, 231, 231, 232, 232, 231, 231, 231, 232, 233, 231, 231, 231, 231, 232, 232, 233, 232, 232, 233, 234, 233, 233, 233, 233, 235, 235, 235, 235, 235, 236, 237, 235, 229, 207, 152, 120, 140, 172, 183, 181, 176, 172, 177, 168, 116, 205, 90, 57, 65, 79, 104, 98, 94, 89, 87, 80, 76, 77, 75, 72, 73, 73, 73, 76, 73, 66, 65, 68, 75, 77, 83, 67, 77, 75, 69, 78, 117, 193, 216, 222, 228, 228, 230, 232, 234, 232, 225, 202, 106, 65, 54, 131, 135, 68, 72, 144, 210, 227, 229, 228, 229, 230, 230, 230, 229, 228, 228, 228, 228, 227, 225, 225, 225, 225, 227, 224, 223, 221, 226, 226, 226, 226, 226, 225, 224, 223, 223, 224, 224, 222, 222, 222, 221, 223, 220, 212, 233, 229, 228, 229, 128, 222, 233, 234, 234, 235, 236, 235, 232, 221, 159, 81, 78, 77, 109, 131, 180, 149, 173, 178, 214, 203, 208, 197, 177, 104, 126, 132, 150, 92, 89, 91, 86, 83, 93, 93, 92, 87, 85, 81, 78, 78, 77, 129, 94, 92, 129, 195, 163, 172, 182, 204, 228, 230, 230, 229, 230, 231, 232, 230, 229, 230, 231, 231, 229, 214, 187, 184, 175, 200, 196, 183, 166, 127, 178, 182, 166, 150, 146, 151, 160, 154, 143, 164, 131, 154, 113, 126, 226, 229, 231, 231, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 230, 230, 229, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 231, 232, 232, 232, 232, 231, 233, 234, 233, 233, 233, 234, 234, 235, 235, 235, 235, 236, 237, 237, 236, 231, 220, 171, 117, 121, 156, 176, 179, 176, 169, 135, 166, 141, 61, 65, 66, 112, 133, 121, 110, 95, 85, 82, 72, 75, 75, 69, 74, 69, 72, 74, 85, 95, 97, 96, 92, 78, 88, 91, 79, 72, 87, 152, 210, 228, 229, 231, 232, 230, 229, 232, 232, 233, 231, 223, 193, 93, 54, 67, 158, 122, 70, 90, 181, 223, 229, 228, 230, 230, 229, 230, 229, 227, 228, 229, 229, 228, 227, 226, 228, 228, 227, 226, 224, 224, 227, 227, 225, 227, 227, 224, 227, 224, 223, 224, 221, 222, 221, 220, 216, 216, 210, 204, 233, 229, 228, 229, 127, 224, 232, 235, 235, 233, 235, 234, 231, 220, 164, 77, 74, 88, 138, 166, 198, 172, 188, 181, 213, 213, 215, 200, 173, 113, 125, 148, 127, 84, 78, 77, 81, 85, 89, 88, 92, 91, 85, 80, 82, 75, 80, 152, 100, 92, 148, 200, 157, 171, 187, 205, 230, 231, 230, 230, 230, 231, 230, 230, 230, 230, 230, 231, 229, 218, 176, 175, 178, 191, 189, 176, 174, 184, 203, 194, 172, 157, 161, 160, 167, 161, 143, 176, 134, 163, 113, 123, 225, 230, 230, 230, 230, 229, 229, 230, 231, 231, 230, 230, 230, 231, 231, 231, 230, 229, 230, 231, 231, 230, 229, 229, 231, 231, 231, 230, 230, 230, 232, 232, 231, 230, 231, 232, 232, 232, 231, 230, 231, 232, 233, 232, 231, 232, 233, 234, 233, 231, 232, 233, 234, 233, 232, 233, 234, 235, 237, 237, 237, 236, 233, 226, 192, 127, 108, 127, 157, 170, 178, 138, 209, 84, 48, 53, 74, 134, 144, 141, 139, 125, 125, 111, 103, 103, 97, 98, 101, 106, 118, 120, 118, 107, 97, 87, 90, 90, 85, 76, 78, 105, 181, 220, 229, 230, 230, 230, 231, 231, 229, 230, 231, 233, 234, 231, 220, 194, 91, 58, 108, 172, 124, 70, 125, 206, 227, 228, 229, 230, 229, 230, 230, 228, 229, 229, 227, 229, 228, 228, 229, 229, 228, 228, 226, 226, 225, 228, 226, 223, 222, 219, 218, 208, 203, 198, 189, 187, 176, 171, 162, 153, 143, 137, 233, 229, 229, 228, 132, 224, 233, 234, 235, 234, 234, 234, 230, 222, 162, 80, 77, 85, 154, 172, 195, 182, 186, 188, 212, 215, 215, 203, 179, 115, 130, 154, 81, 64, 72, 82, 84, 88, 90, 90, 92, 90, 86, 78, 65, 57, 61, 143, 102, 94, 144, 200, 165, 174, 190, 205, 230, 232, 230, 230, 229, 231, 231, 231, 229, 229, 229, 232, 229, 217, 181, 162, 157, 166, 168, 146, 178, 216, 209, 200, 177, 161, 155, 158, 161, 160, 144, 170, 134, 164, 114, 120, 224, 229, 231, 231, 231, 229, 229, 230, 231, 230, 230, 230, 230, 231, 231, 231, 230, 230, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 230, 231, 232, 232, 232, 231, 231, 231, 232, 232, 231, 230, 231, 232, 232, 233, 231, 231, 233, 234, 233, 232, 233, 232, 233, 233, 231, 233, 234, 236, 236, 237, 236, 237, 238, 237, 232, 211, 151, 105, 96, 123, 135, 185, 171, 40, 36, 42, 92, 130, 135, 142, 146, 145, 146, 138, 136, 136, 131, 131, 129, 123, 120, 106, 95, 96, 99, 98, 83, 74, 72, 98, 158, 199, 225, 230, 229, 230, 230, 231, 231, 230, 229, 230, 231, 231, 233, 233, 228, 220, 193, 92, 62, 163, 182, 124, 74, 161, 216, 227, 229, 228, 228, 229, 228, 228, 227, 226, 222, 222, 219, 215, 216, 206, 201, 200, 191, 185, 174, 172, 166, 160, 153, 141, 142, 133, 131, 126, 129, 128, 128, 116, 106, 98, 71, 59, 232, 228, 228, 228, 144, 226, 233, 234, 234, 234, 234, 233, 231, 223, 159, 93, 89, 98, 158, 172, 185, 190, 178, 190, 201, 215, 212, 201, 197, 118, 121, 143, 71, 66, 74, 85, 74, 99, 97, 95, 93, 93, 86, 56, 54, 50, 50, 136, 107, 100, 151, 206, 158, 178, 200, 206, 231, 231, 230, 230, 230, 231, 232, 232, 231, 230, 229, 232, 229, 220, 196, 156, 156, 153, 150, 166, 220, 230, 218, 208, 193, 165, 139, 133, 138, 144, 147, 165, 133, 162, 111, 122, 224, 230, 231, 231, 230, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 231, 232, 230, 230, 230, 232, 232, 231, 231, 231, 231, 232, 231, 231, 231, 230, 232, 233, 232, 231, 231, 232, 233, 233, 232, 232, 232, 234, 234, 234, 233, 234, 234, 236, 236, 236, 236, 237, 239, 239, 235, 225, 189, 131, 112, 140, 209, 76, 40, 39, 46, 109, 137, 136, 126, 125, 124, 119, 114, 117, 114, 104, 102, 98, 99, 96, 109, 102, 93, 84, 57, 56, 77, 122, 184, 212, 223, 226, 226, 227, 227, 227, 227, 229, 227, 226, 225, 226, 228, 229, 230, 230, 224, 215, 189, 72, 136, 198, 158, 99, 107, 177, 197, 194, 190, 185, 179, 177, 169, 161, 162, 154, 144, 144, 134, 135, 131, 126, 126, 126, 118, 117, 121, 122, 124, 123, 117, 122, 113, 101, 89, 79, 64, 55, 46, 42, 43, 53, 52, 233, 229, 229, 230, 135, 226, 233, 234, 234, 234, 234, 235, 230, 222, 155, 92, 91, 88, 159, 165, 176, 201, 177, 191, 189, 214, 211, 207, 199, 131, 148, 105, 67, 72, 72, 76, 87, 99, 98, 96, 96, 87, 62, 44, 48, 51, 48, 132, 100, 102, 152, 200, 158, 181, 199, 208, 230, 230, 230, 230, 229, 231, 232, 232, 231, 229, 229, 228, 227, 222, 206, 180, 167, 157, 185, 222, 232, 232, 230, 213, 205, 180, 157, 159, 157, 155, 164, 160, 134, 163, 111, 120, 225, 230, 231, 231, 230, 230, 230, 230, 231, 231, 231, 230, 230, 231, 231, 231, 230, 230, 230, 232, 231, 231, 230, 230, 231, 231, 232, 231, 230, 230, 232, 232, 232, 231, 231, 231, 232, 232, 231, 231, 231, 232, 233, 232, 231, 231, 232, 233, 233, 232, 231, 232, 233, 234, 234, 233, 233, 234, 235, 236, 235, 236, 237, 238, 239, 240, 237, 235, 226, 187, 185, 175, 50, 34, 35, 46, 106, 137, 141, 138, 140, 147, 139, 136, 131, 111, 124, 109, 121, 112, 100, 89, 57, 45, 39, 38, 40, 52, 64, 91, 114, 125, 137, 148, 153, 156, 157, 155, 155, 153, 147, 154, 152, 153, 148, 155, 153, 148, 127, 109, 68, 80, 94, 89, 94, 95, 107, 112, 110, 115, 109, 119, 106, 106, 108, 113, 120, 115, 116, 118, 116, 118, 112, 113, 116, 117, 112, 102, 88, 79, 74, 60, 54, 43, 41, 42, 44, 50, 67, 79, 94, 100, 106, 112, 233, 230, 230, 232, 147, 227, 234, 232, 233, 234, 235, 235, 231, 221, 143, 78, 75, 89, 159, 164, 175, 198, 176, 193, 185, 214, 211, 203, 203, 136, 159, 74, 65, 74, 68, 77, 93, 99, 95, 103, 94, 81, 47, 46, 46, 45, 47, 138, 103, 96, 147, 197, 156, 189, 205, 212, 230, 230, 230, 229, 230, 230, 231, 230, 229, 229, 229, 229, 230, 225, 215, 219, 219, 212, 225, 230, 232, 233, 233, 226, 216, 197, 165, 152, 157, 147, 155, 160, 134, 170, 113, 135, 227, 230, 231, 232, 231, 230, 229, 230, 231, 231, 231, 230, 230, 231, 231, 230, 229, 230, 230, 231, 231, 231, 230, 230, 231, 232, 231, 230, 231, 231, 232, 232, 232, 231, 231, 232, 232, 232, 232, 232, 232, 233, 232, 232, 231, 232, 232, 233, 233, 232, 232, 232, 233, 234, 234, 233, 234, 234, 235, 236, 234, 236, 236, 239, 238, 239, 237, 238, 236, 184, 222, 112, 170, 136, 79, 46, 43, 56, 69, 85, 91, 110, 109, 107, 98, 89, 95, 66, 65, 52, 48, 50, 49, 52, 50, 48, 49, 50, 54, 56, 59, 59, 67, 68, 78, 74, 74, 78, 77, 79, 76, 72, 73, 75, 77, 78, 78, 73, 67, 64, 60, 62, 71, 72, 72, 73, 77, 82, 86, 91, 97, 102, 105, 106, 103, 101, 105, 107, 100, 96, 87, 85, 69, 63, 56, 48, 46, 43, 51, 45, 43, 49, 60, 73, 77, 90, 100, 116, 121, 125, 130, 128, 124, 117, 233, 229, 229, 232, 154, 229, 234, 233, 235, 235, 236, 236, 232, 221, 138, 79, 75, 85, 153, 156, 165, 181, 165, 175, 167, 199, 188, 183, 183, 135, 139, 70, 66, 70, 78, 77, 95, 97, 98, 106, 97, 67, 47, 42, 44, 49, 45, 145, 105, 97, 161, 205, 166, 189, 195, 211, 230, 231, 229, 229, 230, 231, 230, 230, 229, 230, 230, 228, 228, 219, 211, 219, 214, 210, 215, 215, 231, 233, 233, 231, 224, 209, 184, 163, 164, 156, 154, 156, 133, 174, 118, 132, 226, 230, 232, 231, 230, 230, 230, 230, 230, 231, 231, 230, 230, 231, 231, 230, 230, 230, 230, 232, 231, 231, 230, 230, 231, 231, 232, 231, 231, 231, 232, 232, 231, 231, 231, 232, 233, 232, 232, 232, 232, 234, 233, 232, 230, 219, 218, 231, 233, 230, 232, 233, 234, 234, 235, 234, 234, 234, 235, 233, 231, 229, 225, 224, 216, 206, 200, 191, 187, 196, 163, 77, 113, 99, 64, 44, 47, 49, 52, 53, 55, 57, 59, 54, 52, 50, 51, 51, 52, 48, 51, 55, 51, 57, 53, 54, 48, 53, 49, 51, 52, 52, 60, 56, 62, 60, 57, 57, 63, 57, 59, 58, 59, 64, 58, 60, 58, 53, 53, 59, 60, 58, 64, 66, 75, 74, 77, 74, 78, 76, 76, 73, 79, 70, 62, 58, 51, 48, 44, 46, 44, 46, 48, 48, 51, 57, 61, 82, 81, 88, 98, 109, 106, 109, 111, 121, 119, 129, 128, 132, 131, 118, 110, 98, 234, 232, 230, 234, 147, 232, 236, 237, 236, 238, 239, 239, 235, 225, 137, 82, 74, 83, 99, 91, 100, 94, 93, 99, 116, 131, 122, 114, 121, 144, 94, 77, 90, 91, 79, 82, 78, 65, 72, 109, 101, 57, 50, 52, 57, 53, 50, 146, 107, 106, 168, 211, 160, 190, 196, 208, 230, 231, 230, 228, 230, 231, 230, 230, 229, 229, 230, 229, 229, 211, 200, 210, 199, 208, 209, 205, 222, 232, 233, 233, 229, 220, 208, 186, 190, 180, 154, 149, 135, 178, 113, 139, 227, 230, 232, 232, 231, 230, 230, 231, 232, 231, 230, 230, 230, 231, 231, 231, 231, 230, 231, 232, 232, 231, 231, 231, 231, 232, 233, 231, 232, 232, 233, 233, 233, 232, 232, 234, 234, 234, 233, 234, 235, 237, 237, 232, 226, 212, 136, 195, 194, 174, 202, 211, 214, 211, 210, 203, 192, 189, 182, 164, 151, 133, 124, 112, 98, 89, 80, 80, 90, 156, 66, 60, 54, 50, 53, 49, 55, 54, 55, 55, 58, 57, 51, 54, 50, 57, 55, 58, 54, 56, 53, 58, 56, 53, 57, 45, 53, 50, 49, 51, 50, 53, 48, 53, 59, 57, 54, 53, 49, 54, 52, 55, 55, 58, 55, 53, 53, 50, 58, 64, 94, 94, 84, 68, 69, 72, 66, 53, 51, 49, 45, 41, 38, 40, 41, 49, 61, 75, 73, 80, 93, 100, 111, 104, 116, 117, 118, 120, 129, 130, 132, 130, 130, 129, 119, 123, 117, 120, 115, 122, 121, 110, 104, 101, 235, 232, 230, 235, 139, 231, 237, 237, 236, 239, 240, 240, 235, 226, 133, 90, 73, 77, 64, 65, 66, 66, 71, 74, 95, 99, 119, 140, 153, 158, 71, 78, 94, 82, 68, 63, 52, 54, 52, 91, 103, 56, 72, 97, 103, 70, 51, 140, 98, 107, 168, 207, 157, 184, 189, 215, 231, 230, 230, 228, 231, 231, 231, 230, 230, 231, 230, 230, 228, 218, 205, 201, 196, 196, 201, 199, 213, 232, 233, 233, 231, 228, 221, 220, 225, 216, 173, 143, 137, 178, 109, 138, 226, 230, 232, 233, 231, 230, 230, 231, 231, 232, 231, 231, 231, 232, 233, 232, 231, 231, 231, 233, 232, 232, 232, 232, 231, 234, 234, 233, 233, 234, 235, 235, 235, 234, 235, 236, 237, 238, 237, 238, 240, 242, 244, 240, 234, 222, 114, 85, 79, 86, 86, 82, 80, 84, 89, 86, 84, 86, 78, 79, 75, 72, 67, 70, 66, 69, 64, 67, 62, 66, 55, 56, 58, 58, 64, 64, 62, 63, 91, 95, 60, 51, 51, 53, 47, 56, 51, 50, 53, 51, 81, 62, 77, 54, 63, 54, 59, 53, 53, 52, 51, 51, 53, 54, 82, 64, 67, 57, 51, 52, 47, 55, 49, 52, 50, 49, 52, 46, 57, 76, 128, 85, 72, 53, 47, 41, 40, 40, 35, 50, 58, 67, 81, 96, 96, 116, 127, 131, 132, 136, 149, 142, 145, 138, 137, 131, 127, 121, 128, 127, 119, 122, 124, 123, 115, 115, 115, 107, 109, 113, 115, 106, 111, 108, 234, 231, 230, 235, 135, 230, 237, 237, 238, 238, 240, 239, 235, 226, 126, 95, 78, 77, 55, 60, 64, 68, 71, 85, 109, 165, 210, 220, 216, 167, 77, 77, 71, 68, 60, 53, 53, 54, 51, 74, 121, 64, 99, 120, 119, 80, 58, 135, 99, 106, 171, 211, 152, 188, 191, 216, 231, 231, 230, 230, 230, 230, 231, 230, 230, 231, 231, 231, 229, 222, 214, 196, 186, 191, 192, 185, 205, 232, 233, 234, 232, 232, 227, 225, 226, 219, 168, 146, 132, 176, 109, 136, 225, 230, 232, 232, 232, 231, 231, 232, 232, 233, 231, 232, 231, 232, 233, 232, 231, 231, 232, 232, 233, 232, 232, 232, 228, 233, 235, 233, 233, 234, 234, 235, 235, 235, 235, 237, 238, 238, 239, 240, 241, 244, 245, 241, 232, 214, 85, 72, 64, 65, 64, 61, 60, 62, 58, 84, 71, 75, 56, 59, 54, 58, 57, 57, 51, 53, 72, 54, 60, 53, 48, 50, 48, 48, 52, 56, 58, 78, 102, 106, 55, 53, 49, 48, 49, 48, 46, 51, 49, 47, 104, 67, 69, 50, 50, 49, 45, 50, 50, 48, 51, 49, 54, 70, 111, 80, 62, 48, 48, 46, 52, 54, 52, 50, 50, 49, 44, 46, 56, 65, 98, 64, 85, 102, 91, 82, 81, 82, 95, 101, 119, 135, 144, 148, 144, 153, 145, 141, 131, 126, 129, 129, 127, 129, 127, 121, 126, 124, 124, 120, 118, 122, 115, 117, 110, 110, 102, 104, 109, 117, 125, 131, 122, 117, 233, 232, 229, 234, 144, 231, 237, 237, 236, 238, 240, 238, 234, 224, 121, 87, 76, 81, 63, 70, 86, 103, 86, 135, 186, 227, 231, 231, 220, 123, 60, 73, 59, 84, 80, 56, 60, 73, 65, 68, 128, 73, 88, 110, 114, 87, 64, 139, 97, 102, 170, 210, 152, 185, 180, 216, 230, 231, 229, 229, 230, 231, 230, 231, 229, 231, 232, 231, 229, 219, 211, 188, 185, 186, 183, 163, 202, 232, 233, 233, 232, 232, 231, 226, 225, 219, 169, 145, 132, 167, 113, 137, 227, 230, 232, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 232, 233, 232, 230, 231, 232, 232, 233, 232, 232, 232, 230, 233, 234, 233, 233, 234, 234, 230, 233, 234, 236, 238, 239, 239, 240, 241, 242, 244, 245, 241, 232, 206, 85, 68, 57, 59, 51, 60, 60, 60, 50, 90, 82, 61, 63, 50, 44, 50, 51, 50, 49, 47, 83, 56, 58, 53, 48, 46, 45, 44, 48, 48, 56, 96, 102, 111, 51, 48, 45, 45, 46, 47, 46, 50, 45, 46, 98, 67, 68, 47, 50, 45, 43, 49, 46, 46, 54, 47, 52, 82, 106, 83, 60, 48, 47, 45, 46, 49, 47, 51, 43, 48, 47, 46, 68, 65, 74, 66, 109, 121, 122, 127, 138, 137, 145, 149, 149, 144, 131, 124, 120, 121, 116, 122, 122, 126, 138, 129, 122, 121, 113, 112, 111, 117, 114, 122, 119, 117, 123, 121, 116, 119, 118, 114, 113, 119, 112, 112, 102, 90, 233, 230, 229, 233, 135, 231, 236, 236, 235, 236, 238, 236, 231, 220, 115, 85, 74, 93, 90, 122, 162, 152, 111, 160, 225, 233, 236, 229, 217, 89, 59, 77, 70, 86, 74, 60, 72, 100, 81, 82, 138, 101, 74, 95, 84, 81, 62, 139, 92, 108, 168, 203, 154, 186, 186, 218, 230, 230, 230, 230, 230, 230, 229, 227, 229, 229, 231, 231, 228, 212, 206, 190, 189, 189, 179, 175, 224, 233, 233, 233, 233, 232, 232, 228, 227, 220, 169, 145, 131, 157, 106, 142, 228, 231, 231, 232, 232, 231, 231, 232, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 232, 232, 233, 232, 232, 232, 234, 234, 234, 233, 232, 232, 221, 220, 229, 231, 236, 238, 239, 240, 240, 241, 242, 245, 246, 242, 231, 206, 80, 64, 55, 49, 49, 50, 51, 56, 54, 87, 78, 56, 54, 49, 46, 44, 47, 50, 52, 45, 93, 57, 59, 50, 46, 46, 41, 42, 45, 50, 56, 117, 103, 90, 50, 45, 50, 47, 45, 46, 48, 46, 50, 46, 103, 57, 67, 48, 45, 46, 44, 48, 47, 45, 46, 44, 53, 82, 95, 92, 55, 49, 49, 44, 48, 43, 42, 47, 48, 50, 44, 41, 70, 74, 63, 97, 149, 147, 134, 124, 111, 110, 108, 114, 115, 109, 119, 114, 112, 110, 119, 120, 124, 129, 123, 126, 118, 123, 112, 106, 112, 113, 120, 122, 115, 119, 114, 112, 112, 113, 106, 103, 97, 101, 93, 89, 85, 82, 232, 229, 229, 232, 149, 231, 235, 235, 235, 237, 238, 236, 230, 220, 113, 86, 80, 104, 150, 161, 146, 122, 106, 178, 231, 238, 235, 226, 202, 72, 62, 67, 70, 61, 54, 67, 81, 94, 82, 98, 138, 113, 104, 85, 86, 70, 62, 141, 85, 118, 158, 177, 155, 190, 179, 216, 230, 230, 230, 230, 229, 230, 229, 229, 230, 231, 230, 228, 227, 195, 199, 188, 188, 185, 180, 215, 230, 232, 233, 233, 232, 232, 232, 227, 227, 220, 197, 147, 131, 177, 108, 142, 228, 231, 232, 232, 231, 231, 231, 232, 233, 232, 232, 231, 231, 232, 232, 232, 230, 231, 232, 233, 233, 233, 233, 232, 234, 234, 227, 232, 234, 231, 232, 236, 231, 234, 232, 238, 239, 240, 240, 236, 243, 245, 246, 243, 230, 201, 71, 56, 56, 62, 53, 51, 52, 53, 50, 98, 76, 48, 46, 52, 46, 47, 46, 49, 51, 46, 73, 56, 56, 49, 45, 48, 44, 42, 48, 49, 50, 91, 91, 80, 49, 46, 48, 42, 46, 46, 48, 47, 53, 45, 113, 71, 72, 70, 46, 46, 48, 50, 48, 40, 47, 47, 60, 108, 94, 107, 61, 51, 45, 43, 46, 52, 45, 46, 53, 47, 48, 53, 85, 83, 57, 90, 110, 103, 97, 95, 103, 97, 101, 106, 107, 112, 110, 114, 115, 116, 122, 112, 113, 124, 123, 122, 121, 114, 112, 112, 110, 114, 116, 112, 109, 109, 112, 106, 104, 100, 89, 81, 80, 92, 83, 91, 87, 83, 233, 230, 230, 233, 137, 230, 234, 235, 235, 236, 237, 235, 230, 220, 105, 86, 81, 111, 146, 149, 135, 115, 163, 214, 232, 237, 237, 227, 205, 75, 60, 59, 58, 75, 56, 60, 82, 73, 77, 99, 138, 97, 107, 87, 118, 91, 60, 135, 80, 124, 169, 182, 149, 187, 167, 219, 229, 230, 229, 229, 230, 230, 230, 229, 229, 230, 231, 228, 227, 204, 192, 185, 184, 183, 188, 227, 231, 232, 233, 233, 231, 232, 233, 232, 229, 223, 208, 148, 130, 173, 107, 136, 227, 230, 231, 232, 231, 230, 231, 230, 233, 232, 232, 231, 231, 233, 232, 231, 231, 231, 232, 233, 233, 232, 232, 232, 234, 234, 228, 231, 233, 234, 235, 236, 236, 236, 236, 238, 239, 240, 239, 240, 242, 245, 246, 242, 230, 191, 71, 59, 59, 51, 55, 55, 43, 63, 48, 79, 81, 50, 49, 53, 48, 50, 50, 52, 52, 47, 81, 58, 51, 45, 45, 48, 42, 46, 42, 49, 50, 82, 80, 69, 51, 45, 50, 46, 48, 52, 47, 53, 52, 46, 105, 69, 66, 88, 57, 54, 56, 54, 57, 47, 93, 57, 65, 131, 99, 105, 52, 47, 49, 45, 50, 45, 46, 49, 46, 52, 50, 53, 95, 94, 58, 70, 102, 95, 96, 101, 96, 100, 97, 104, 113, 107, 114, 111, 112, 112, 106, 107, 108, 111, 111, 109, 110, 105, 96, 99, 101, 103, 106, 97, 100, 104, 104, 98, 87, 84, 82, 80, 89, 105, 97, 100, 98, 88, 233, 230, 230, 234, 144, 230, 235, 234, 234, 235, 235, 233, 227, 218, 102, 85, 83, 115, 171, 188, 160, 188, 216, 227, 233, 237, 236, 226, 197, 74, 56, 54, 64, 69, 78, 75, 95, 95, 94, 98, 148, 79, 92, 88, 103, 88, 61, 136, 83, 115, 173, 182, 144, 177, 161, 216, 227, 229, 230, 230, 230, 230, 229, 226, 228, 230, 231, 230, 228, 216, 184, 180, 174, 175, 200, 230, 231, 232, 233, 233, 232, 232, 233, 233, 230, 223, 208, 155, 128, 173, 110, 134, 227, 230, 231, 232, 231, 231, 231, 232, 232, 232, 232, 230, 231, 232, 233, 232, 231, 231, 232, 233, 234, 232, 232, 232, 234, 234, 231, 227, 234, 235, 236, 236, 236, 236, 237, 238, 239, 240, 240, 241, 242, 245, 245, 242, 230, 181, 77, 53, 57, 55, 53, 48, 48, 53, 48, 71, 87, 49, 49, 51, 48, 51, 51, 45, 52, 46, 67, 57, 51, 47, 45, 45, 46, 48, 46, 47, 50, 72, 64, 66, 50, 45, 48, 43, 46, 49, 44, 50, 57, 49, 110, 70, 68, 81, 78, 91, 96, 95, 99, 57, 84, 99, 66, 137, 93, 103, 52, 50, 47, 45, 44, 44, 47, 45, 48, 47, 50, 62, 86, 96, 55, 84, 103, 95, 100, 102, 107, 101, 101, 107, 105, 103, 103, 103, 103, 97, 95, 102, 101, 99, 102, 107, 104, 100, 93, 90, 89, 92, 96, 97, 96, 99, 103, 106, 98, 95, 96, 97, 90, 107, 101, 96, 102, 96, 232, 229, 229, 234, 137, 229, 234, 234, 234, 234, 235, 233, 227, 215, 94, 87, 82, 113, 149, 203, 206, 213, 219, 231, 235, 235, 234, 228, 163, 134, 59, 53, 62, 88, 125, 80, 97, 98, 80, 104, 146, 88, 93, 73, 78, 78, 72, 145, 84, 122, 172, 183, 144, 183, 170, 218, 228, 229, 228, 229, 230, 230, 229, 227, 229, 230, 231, 229, 225, 211, 175, 168, 162, 165, 216, 230, 232, 232, 232, 233, 232, 232, 232, 234, 231, 222, 208, 161, 131, 178, 114, 135, 226, 230, 231, 232, 231, 231, 231, 231, 233, 233, 231, 231, 231, 232, 233, 233, 232, 231, 231, 233, 233, 233, 232, 233, 234, 235, 234, 234, 234, 234, 236, 235, 236, 236, 237, 238, 240, 241, 240, 241, 242, 245, 246, 242, 230, 172, 71, 56, 56, 56, 48, 46, 48, 54, 52, 84, 78, 54, 49, 49, 51, 52, 47, 51, 49, 48, 73, 63, 53, 50, 44, 47, 47, 48, 45, 51, 51, 78, 67, 75, 50, 54, 50, 42, 47, 43, 48, 47, 52, 49, 108, 76, 74, 68, 88, 73, 76, 81, 90, 55, 86, 76, 67, 128, 81, 112, 52, 46, 45, 44, 41, 40, 44, 43, 48, 46, 49, 69, 86, 108, 47, 111, 101, 106, 101, 97, 93, 99, 98, 100, 100, 94, 99, 93, 99, 102, 107, 104, 110, 108, 110, 117, 115, 113, 106, 105, 102, 105, 106, 102, 98, 103, 102, 100, 97, 91, 90, 90, 91, 111, 114, 114, 121, 100, 233, 229, 229, 232, 132, 228, 233, 234, 233, 233, 235, 231, 226, 213, 94, 90, 87, 116, 189, 207, 211, 215, 220, 230, 234, 231, 228, 220, 92, 155, 122, 60, 108, 142, 146, 126, 91, 92, 80, 144, 150, 107, 84, 79, 73, 76, 106, 149, 77, 110, 178, 180, 148, 192, 166, 219, 228, 230, 228, 229, 230, 229, 229, 230, 229, 231, 230, 228, 223, 194, 163, 157, 160, 183, 225, 230, 231, 232, 233, 233, 232, 232, 232, 233, 230, 222, 203, 163, 131, 175, 108, 135, 227, 230, 232, 232, 232, 231, 231, 231, 232, 232, 231, 231, 231, 232, 233, 232, 231, 230, 231, 232, 233, 232, 232, 232, 234, 235, 234, 233, 234, 235, 236, 236, 236, 236, 237, 238, 240, 240, 240, 241, 241, 245, 246, 242, 230, 171, 72, 59, 54, 50, 54, 51, 55, 56, 56, 90, 76, 52, 48, 46, 47, 46, 48, 53, 50, 49, 81, 64, 54, 46, 47, 46, 45, 49, 49, 50, 54, 76, 62, 64, 52, 57, 48, 46, 42, 48, 45, 47, 50, 52, 99, 77, 70, 77, 83, 81, 66, 79, 75, 58, 91, 80, 64, 136, 77, 117, 53, 43, 48, 49, 45, 42, 45, 44, 40, 50, 51, 92, 89, 112, 49, 91, 92, 93, 96, 96, 94, 89, 93, 93, 95, 94, 96, 106, 111, 110, 111, 110, 112, 115, 121, 114, 115, 116, 110, 108, 103, 102, 111, 100, 102, 108, 112, 106, 105, 105, 105, 106, 111, 116, 117, 104, 110, 110, 230, 229, 228, 232, 136, 229, 233, 234, 233, 234, 235, 233, 225, 211, 94, 91, 92, 125, 201, 214, 215, 221, 225, 228, 233, 231, 225, 204, 102, 108, 160, 105, 147, 158, 158, 155, 135, 125, 104, 166, 149, 113, 62, 71, 75, 93, 172, 141, 76, 110, 179, 174, 146, 190, 170, 222, 228, 230, 229, 229, 230, 230, 231, 230, 230, 231, 229, 225, 212, 176, 157, 152, 152, 199, 230, 230, 231, 232, 232, 233, 232, 232, 233, 233, 230, 224, 201, 153, 131, 171, 106, 139, 227, 231, 231, 233, 232, 231, 231, 231, 232, 233, 232, 231, 231, 233, 233, 232, 231, 231, 232, 233, 233, 232, 232, 232, 234, 234, 234, 233, 234, 234, 236, 236, 236, 236, 236, 238, 240, 240, 240, 241, 242, 245, 245, 241, 229, 166, 70, 57, 53, 67, 58, 60, 57, 58, 57, 89, 78, 49, 47, 52, 45, 50, 46, 49, 51, 53, 90, 65, 48, 45, 46, 45, 42, 48, 48, 53, 51, 77, 63, 70, 51, 47, 44, 50, 44, 46, 41, 44, 52, 54, 106, 80, 70, 84, 81, 95, 59, 63, 55, 59, 92, 75, 57, 126, 85, 113, 49, 48, 48, 46, 43, 42, 41, 44, 47, 47, 52, 96, 83, 115, 45, 73, 83, 91, 102, 99, 93, 93, 99, 108, 105, 108, 102, 108, 113, 106, 115, 112, 113, 118, 126, 122, 119, 120, 114, 113, 114, 112, 111, 106, 112, 108, 112, 112, 112, 100, 99, 100, 103, 108, 113, 107, 108, 117, 231, 229, 229, 231, 151, 228, 232, 234, 233, 233, 235, 233, 223, 210, 94, 88, 98, 128, 204, 216, 218, 218, 222, 224, 227, 231, 225, 196, 147, 103, 152, 127, 156, 176, 189, 170, 166, 161, 154, 146, 137, 73, 61, 70, 92, 146, 191, 131, 82, 133, 172, 173, 146, 187, 161, 220, 228, 230, 229, 228, 230, 231, 230, 230, 228, 227, 220, 213, 193, 169, 155, 148, 154, 209, 225, 229, 230, 230, 231, 231, 230, 231, 232, 233, 230, 223, 203, 147, 131, 169, 107, 138, 227, 230, 231, 229, 231, 231, 231, 231, 232, 233, 231, 231, 231, 232, 232, 232, 231, 231, 232, 233, 233, 232, 232, 232, 234, 234, 234, 233, 233, 235, 236, 236, 236, 236, 236, 238, 240, 240, 240, 241, 242, 245, 245, 240, 228, 178, 65, 56, 67, 62, 59, 63, 64, 57, 59, 105, 73, 46, 60, 49, 42, 70, 46, 50, 48, 43, 83, 64, 49, 47, 48, 46, 47, 47, 47, 46, 53, 88, 71, 74, 49, 44, 48, 45, 46, 46, 44, 46, 55, 58, 104, 78, 65, 69, 50, 60, 125, 58, 49, 54, 90, 81, 57, 139, 87, 118, 51, 45, 50, 47, 46, 38, 41, 49, 49, 41, 48, 100, 85, 118, 58, 91, 98, 94, 94, 100, 101, 101, 97, 94, 95, 91, 100, 101, 114, 111, 112, 110, 119, 119, 121, 120, 126, 117, 116, 113, 110, 106, 108, 105, 113, 109, 107, 106, 107, 102, 99, 97, 103, 107, 109, 112, 118, 120, 232, 228, 229, 233, 146, 229, 233, 234, 233, 234, 235, 233, 224, 209, 92, 88, 101, 128, 205, 212, 214, 218, 218, 221, 223, 228, 225, 181, 147, 140, 135, 107, 162, 210, 213, 199, 170, 160, 152, 147, 99, 68, 93, 90, 115, 191, 192, 129, 84, 130, 184, 190, 149, 190, 162, 222, 231, 230, 229, 229, 229, 230, 228, 226, 219, 211, 200, 186, 174, 161, 149, 134, 176, 204, 206, 203, 198, 194, 205, 206, 206, 212, 215, 227, 230, 222, 203, 158, 125, 172, 105, 146, 228, 230, 231, 231, 232, 231, 231, 232, 233, 232, 231, 232, 231, 232, 232, 232, 231, 231, 232, 233, 233, 232, 232, 233, 234, 234, 234, 233, 234, 234, 236, 236, 236, 236, 236, 238, 239, 240, 240, 240, 242, 245, 245, 242, 230, 191, 75, 58, 84, 61, 58, 60, 58, 63, 60, 99, 72, 48, 51, 50, 44, 48, 46, 45, 50, 42, 75, 65, 47, 44, 44, 51, 46, 51, 47, 46, 48, 76, 66, 74, 49, 47, 44, 40, 40, 42, 41, 46, 49, 52, 99, 74, 65, 72, 80, 77, 106, 71, 55, 53, 86, 85, 90, 157, 97, 114, 46, 43, 43, 45, 53, 41, 43, 43, 47, 48, 48, 96, 87, 109, 60, 82, 101, 93, 106, 104, 110, 106, 102, 101, 106, 98, 104, 106, 110, 117, 117, 117, 121, 124, 122, 126, 123, 119, 120, 113, 105, 108, 103, 104, 104, 105, 106, 109, 111, 109, 109, 109, 110, 114, 118, 121, 111, 110, 233, 228, 228, 231, 138, 228, 233, 234, 234, 234, 235, 232, 223, 206, 85, 88, 100, 129, 203, 216, 215, 207, 195, 201, 209, 219, 217, 122, 108, 146, 142, 100, 181, 216, 213, 206, 169, 148, 144, 146, 126, 136, 116, 102, 169, 199, 190, 130, 85, 143, 186, 182, 139, 192, 161, 223, 231, 232, 230, 226, 225, 221, 210, 206, 195, 183, 172, 168, 162, 137, 128, 126, 194, 166, 128, 146, 168, 181, 197, 200, 198, 195, 202, 210, 227, 222, 203, 166, 136, 173, 113, 139, 228, 230, 232, 232, 232, 231, 231, 232, 232, 233, 232, 231, 232, 232, 232, 231, 232, 231, 232, 233, 233, 232, 232, 232, 233, 234, 234, 233, 233, 234, 236, 235, 235, 236, 236, 238, 239, 239, 239, 240, 242, 243, 245, 241, 229, 203, 75, 65, 127, 64, 73, 64, 65, 65, 55, 93, 74, 52, 48, 44, 47, 42, 42, 51, 49, 46, 79, 67, 48, 47, 46, 47, 47, 44, 45, 46, 51, 77, 69, 75, 52, 46, 46, 43, 42, 44, 44, 44, 49, 59, 109, 69, 68, 66, 49, 67, 105, 101, 89, 57, 86, 88, 53, 144, 86, 100, 48, 48, 45, 48, 41, 43, 42, 40, 42, 54, 54, 116, 91, 91, 55, 92, 105, 97, 100, 112, 105, 96, 102, 103, 102, 103, 104, 119, 112, 113, 119, 117, 122, 122, 120, 128, 126, 122, 122, 115, 110, 107, 99, 101, 108, 107, 107, 111, 107, 118, 114, 118, 120, 117, 107, 101, 93, 100, 234, 231, 229, 231, 129, 226, 234, 235, 234, 235, 236, 233, 224, 204, 92, 83, 105, 127, 207, 215, 210, 198, 147, 120, 160, 195, 206, 67, 49, 93, 132, 121, 194, 218, 218, 197, 165, 142, 116, 128, 143, 170, 125, 144, 205, 206, 197, 133, 89, 140, 192, 183, 149, 190, 161, 225, 230, 229, 224, 222, 202, 193, 180, 177, 168, 160, 146, 132, 122, 109, 108, 116, 127, 123, 122, 140, 157, 169, 201, 194, 190, 197, 202, 208, 227, 223, 205, 166, 137, 179, 115, 140, 228, 230, 232, 232, 232, 231, 231, 231, 232, 232, 231, 231, 231, 232, 232, 233, 231, 231, 232, 233, 233, 232, 232, 232, 233, 234, 234, 233, 233, 234, 235, 236, 235, 235, 236, 238, 239, 239, 239, 240, 242, 244, 245, 241, 230, 209, 84, 64, 149, 66, 62, 64, 65, 65, 54, 101, 65, 43, 45, 48, 45, 42, 46, 43, 52, 45, 76, 62, 50, 45, 45, 48, 48, 45, 48, 48, 48, 80, 72, 74, 46, 46, 48, 46, 42, 42, 41, 46, 49, 60, 115, 78, 65, 71, 62, 63, 109, 78, 54, 50, 94, 95, 58, 145, 80, 93, 44, 46, 44, 42, 39, 40, 42, 39, 45, 42, 47, 110, 89, 104, 67, 85, 89, 94, 97, 105, 101, 105, 105, 105, 110, 109, 111, 112, 112, 113, 112, 121, 121, 118, 117, 126, 122, 120, 120, 112, 112, 110, 100, 105, 103, 105, 108, 106, 101, 111, 98, 95, 93, 97, 92, 98, 96, 92, 234, 231, 229, 232, 139, 228, 234, 235, 235, 235, 236, 234, 225, 201, 95, 85, 108, 126, 205, 216, 205, 192, 129, 128, 145, 181, 187, 51, 54, 54, 111, 132, 183, 212, 197, 182, 113, 98, 84, 101, 150, 150, 129, 196, 214, 208, 197, 125, 86, 148, 199, 181, 154, 190, 166, 223, 227, 218, 214, 192, 176, 170, 158, 140, 119, 117, 98, 90, 86, 88, 100, 103, 100, 108, 117, 137, 148, 160, 170, 181, 187, 192, 198, 209, 224, 222, 204, 162, 137, 181, 111, 138, 228, 230, 232, 231, 232, 231, 231, 231, 232, 232, 231, 231, 231, 233, 233, 233, 232, 232, 232, 233, 233, 232, 232, 232, 232, 234, 234, 233, 233, 234, 235, 236, 235, 235, 236, 238, 239, 239, 239, 241, 242, 244, 245, 241, 230, 213, 81, 62, 157, 64, 63, 65, 72, 64, 51, 95, 76, 50, 48, 44, 42, 45, 44, 46, 46, 43, 80, 59, 50, 45, 47, 49, 46, 45, 41, 47, 53, 71, 67, 69, 48, 42, 45, 45, 39, 44, 41, 45, 54, 55, 123, 72, 66, 69, 65, 62, 58, 46, 50, 46, 53, 93, 60, 147, 73, 92, 47, 46, 46, 40, 42, 43, 42, 43, 47, 43, 51, 118, 96, 102, 69, 79, 85, 90, 98, 98, 105, 111, 107, 108, 109, 108, 111, 109, 113, 119, 111, 103, 113, 110, 115, 117, 110, 112, 116, 112, 107, 110, 106, 101, 101, 96, 103, 100, 90, 90, 88, 97, 92, 104, 106, 104, 106, 104, 234, 231, 228, 231, 120, 225, 235, 235, 235, 236, 237, 235, 225, 204, 89, 88, 106, 121, 194, 193, 169, 160, 122, 119, 132, 153, 170, 67, 80, 81, 78, 129, 155, 122, 105, 104, 87, 75, 85, 121, 158, 148, 152, 217, 217, 211, 195, 125, 92, 143, 201, 174, 156, 196, 170, 216, 222, 216, 194, 150, 128, 114, 100, 98, 93, 87, 80, 84, 89, 107, 103, 117, 108, 110, 128, 141, 153, 163, 175, 180, 185, 189, 197, 207, 227, 223, 205, 165, 128, 181, 109, 134, 227, 230, 231, 231, 232, 231, 230, 231, 232, 232, 231, 231, 231, 232, 233, 233, 232, 232, 232, 233, 233, 233, 232, 233, 233, 234, 234, 233, 233, 234, 235, 236, 236, 236, 236, 237, 239, 240, 240, 241, 242, 244, 245, 242, 232, 219, 82, 53, 121, 60, 66, 63, 62, 62, 47, 89, 57, 47, 42, 45, 48, 45, 49, 47, 56, 42, 82, 61, 55, 45, 44, 45, 41, 43, 43, 48, 49, 77, 72, 73, 50, 47, 49, 41, 43, 39, 45, 51, 49, 49, 114, 70, 64, 71, 64, 59, 70, 60, 78, 48, 85, 48, 51, 129, 72, 91, 51, 43, 43, 47, 41, 41, 40, 41, 47, 44, 46, 94, 95, 89, 81, 88, 88, 91, 97, 106, 109, 115, 121, 116, 113, 108, 111, 115, 112, 113, 109, 105, 109, 111, 108, 113, 113, 112, 107, 98, 94, 90, 94, 96, 102, 96, 105, 95, 97, 93, 95, 97, 109, 108, 114, 116, 106, 102, 234, 232, 231, 233, 150, 230, 235, 237, 236, 238, 239, 237, 227, 207, 91, 84, 100, 108, 167, 102, 80, 96, 103, 107, 119, 137, 160, 110, 82, 59, 60, 132, 144, 84, 91, 97, 83, 74, 105, 130, 151, 136, 183, 216, 213, 203, 194, 115, 92, 145, 179, 144, 155, 199, 180, 218, 217, 206, 172, 153, 157, 170, 171, 172, 166, 145, 131, 129, 135, 142, 146, 152, 152, 135, 142, 147, 167, 187, 185, 185, 184, 187, 189, 207, 226, 224, 209, 171, 129, 176, 106, 141, 228, 230, 231, 231, 232, 231, 231, 231, 232, 232, 231, 231, 230, 232, 232, 233, 232, 232, 232, 233, 234, 233, 232, 233, 234, 234, 234, 233, 233, 234, 235, 236, 236, 236, 236, 238, 239, 240, 240, 241, 242, 244, 246, 242, 234, 220, 82, 51, 67, 73, 67, 80, 64, 56, 48, 91, 56, 47, 50, 49, 44, 47, 45, 47, 48, 47, 80, 61, 54, 47, 45, 45, 46, 50, 45, 43, 49, 70, 73, 75, 48, 47, 45, 42, 42, 45, 41, 48, 47, 48, 119, 70, 62, 73, 56, 62, 89, 91, 90, 56, 87, 61, 54, 124, 82, 90, 53, 46, 43, 48, 41, 40, 38, 43, 46, 47, 52, 83, 100, 97, 66, 97, 124, 122, 118, 108, 103, 98, 101, 99, 98, 93, 92, 101, 100, 111, 108, 98, 106, 110, 113, 117, 114, 109, 102, 96, 91, 95, 98, 99, 102, 105, 107, 102, 104, 105, 104, 108, 108, 110, 112, 108, 98, 85, 235, 232, 231, 233, 136, 229, 237, 238, 238, 239, 240, 238, 228, 206, 92, 81, 97, 105, 145, 78, 87, 86, 98, 107, 104, 116, 107, 45, 41, 44, 46, 131, 147, 95, 67, 73, 96, 90, 143, 157, 173, 181, 208, 220, 213, 198, 189, 107, 92, 157, 190, 143, 144, 201, 163, 218, 219, 195, 157, 170, 193, 196, 203, 203, 206, 189, 162, 167, 168, 170, 178, 175, 173, 173, 160, 170, 165, 186, 177, 164, 167, 174, 192, 204, 225, 227, 220, 176, 125, 185, 109, 141, 228, 231, 231, 231, 232, 231, 231, 231, 232, 232, 232, 232, 231, 231, 232, 232, 232, 232, 232, 234, 234, 233, 232, 232, 233, 234, 234, 234, 234, 235, 235, 236, 236, 236, 237, 238, 239, 240, 240, 241, 242, 244, 246, 243, 236, 225, 95, 57, 55, 63, 56, 60, 62, 52, 46, 93, 59, 51, 46, 41, 42, 50, 41, 45, 50, 47, 74, 59, 55, 51, 48, 52, 50, 46, 47, 46, 52, 58, 73, 77, 50, 49, 48, 43, 39, 44, 46, 48, 46, 44, 108, 64, 70, 84, 58, 69, 52, 51, 62, 44, 71, 85, 65, 104, 79, 80, 49, 42, 43, 42, 44, 39, 40, 43, 40, 46, 51, 80, 98, 108, 56, 112, 130, 117, 115, 105, 100, 93, 96, 96, 98, 103, 97, 102, 106, 112, 105, 111, 105, 110, 112, 108, 112, 109, 100, 107, 97, 103, 105, 105, 103, 107, 107, 105, 94, 95, 93, 90, 103, 101, 99, 110, 104, 94, 235, 231, 232, 234, 143, 231, 237, 238, 239, 239, 239, 237, 228, 201, 90, 78, 97, 88, 117, 82, 99, 91, 86, 82, 89, 108, 80, 37, 38, 48, 47, 141, 164, 134, 103, 116, 143, 176, 209, 210, 195, 197, 209, 218, 213, 202, 186, 111, 102, 164, 201, 140, 155, 209, 174, 220, 220, 182, 182, 166, 189, 189, 196, 197, 204, 190, 164, 163, 168, 175, 170, 177, 176, 177, 175, 158, 163, 145, 148, 168, 166, 174, 186, 200, 225, 227, 222, 186, 126, 178, 109, 136, 228, 231, 231, 231, 231, 231, 231, 231, 232, 233, 232, 231, 231, 232, 233, 233, 232, 232, 232, 234, 233, 232, 233, 232, 233, 234, 235, 234, 234, 234, 236, 236, 236, 236, 237, 238, 240, 239, 240, 241, 242, 244, 246, 244, 238, 227, 111, 48, 52, 44, 52, 57, 53, 43, 43, 102, 62, 52, 47, 44, 47, 46, 45, 47, 49, 48, 67, 55, 56, 46, 41, 41, 42, 47, 46, 44, 48, 58, 74, 76, 51, 47, 48, 46, 42, 40, 42, 50, 42, 45, 103, 62, 75, 87, 62, 62, 53, 61, 52, 47, 69, 66, 55, 97, 83, 87, 46, 43, 47, 41, 45, 39, 42, 42, 44, 42, 51, 64, 94, 100, 50, 94, 89, 100, 101, 96, 103, 103, 100, 103, 104, 99, 99, 99, 98, 108, 105, 108, 106, 108, 112, 111, 113, 111, 110, 107, 104, 107, 99, 97, 98, 106, 107, 103, 98, 95, 92, 93, 105, 100, 102, 114, 107, 98, 234, 232, 232, 235, 158, 232, 237, 238, 238, 239, 239, 237, 228, 198, 90, 74, 87, 75, 88, 85, 97, 102, 85, 98, 87, 112, 61, 32, 38, 42, 45, 152, 167, 164, 154, 142, 158, 172, 202, 216, 194, 203, 211, 220, 218, 202, 187, 104, 99, 162, 206, 145, 153, 207, 156, 217, 217, 166, 178, 143, 160, 167, 166, 171, 182, 184, 153, 160, 161, 162, 164, 167, 165, 166, 166, 155, 153, 143, 144, 155, 157, 170, 179, 197, 221, 227, 224, 202, 131, 184, 110, 142, 229, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 231, 232, 232, 232, 232, 232, 232, 234, 233, 233, 233, 232, 233, 234, 234, 234, 234, 234, 235, 236, 236, 236, 236, 237, 239, 239, 239, 240, 241, 244, 246, 244, 239, 227, 127, 52, 54, 49, 46, 51, 49, 44, 47, 91, 60, 56, 49, 49, 43, 45, 42, 41, 43, 46, 64, 59, 58, 45, 42, 42, 42, 47, 44, 49, 53, 53, 87, 76, 59, 45, 44, 41, 40, 42, 40, 46, 48, 43, 93, 60, 71, 76, 52, 51, 45, 79, 70, 52, 64, 61, 53, 73, 78, 91, 49, 42, 45, 40, 43, 36, 39, 38, 42, 43, 48, 61, 107, 112, 58, 91, 87, 98, 93, 96, 103, 91, 92, 93, 105, 104, 105, 112, 105, 102, 100, 102, 97, 107, 109, 109, 110, 108, 106, 105, 97, 94, 97, 94, 100, 106, 100, 100, 97, 96, 99, 96, 98, 110, 104, 115, 115, 96, 235, 232, 231, 236, 135, 233, 237, 238, 238, 239, 239, 237, 228, 193, 83, 72, 86, 73, 97, 82, 95, 95, 93, 83, 99, 127, 52, 38, 39, 45, 51, 157, 163, 153, 115, 87, 88, 136, 204, 215, 202, 212, 219, 220, 218, 204, 186, 100, 109, 156, 211, 137, 160, 202, 156, 218, 219, 183, 180, 127, 121, 113, 109, 117, 134, 152, 139, 148, 147, 151, 153, 160, 158, 158, 154, 153, 146, 143, 152, 157, 158, 167, 173, 192, 218, 223, 223, 210, 128, 183, 108, 146, 228, 230, 231, 232, 232, 231, 230, 231, 232, 231, 231, 231, 231, 231, 232, 226, 231, 232, 233, 234, 234, 233, 233, 233, 234, 234, 234, 233, 233, 234, 235, 236, 236, 236, 236, 238, 239, 240, 240, 240, 242, 244, 246, 244, 240, 227, 141, 52, 44, 46, 49, 50, 49, 44, 51, 80, 63, 59, 48, 47, 50, 41, 41, 51, 45, 48, 61, 60, 57, 45, 44, 41, 46, 47, 49, 49, 52, 46, 77, 73, 47, 46, 51, 52, 45, 43, 43, 49, 51, 49, 96, 61, 78, 72, 67, 55, 45, 68, 56, 45, 66, 69, 50, 70, 83, 75, 46, 43, 45, 39, 37, 43, 37, 40, 42, 42, 52, 50, 97, 103, 52, 76, 80, 96, 102, 94, 102, 98, 94, 103, 108, 97, 100, 99, 97, 105, 114, 114, 120, 124, 116, 112, 104, 108, 102, 104, 103, 99, 108, 101, 106, 108, 105, 109, 104, 108, 97, 97, 93, 100, 91, 89, 88, 69, 236, 231, 231, 235, 133, 232, 237, 238, 238, 239, 239, 237, 227, 189, 86, 76, 92, 92, 118, 82, 84, 92, 91, 80, 128, 134, 43, 40, 43, 52, 59, 151, 150, 105, 96, 95, 86, 114, 189, 216, 181, 206, 220, 222, 216, 199, 176, 98, 109, 153, 209, 142, 161, 205, 164, 227, 227, 212, 200, 182, 121, 119, 134, 129, 106, 110, 115, 114, 127, 136, 136, 146, 152, 145, 145, 142, 131, 140, 137, 152, 153, 158, 168, 188, 214, 217, 220, 213, 124, 180, 102, 150, 228, 231, 231, 232, 232, 231, 231, 231, 232, 232, 231, 231, 230, 232, 230, 229, 230, 231, 232, 234, 234, 233, 233, 233, 233, 234, 234, 233, 233, 234, 236, 235, 236, 236, 236, 238, 239, 240, 240, 240, 242, 244, 246, 244, 241, 228, 161, 57, 49, 43, 46, 50, 43, 45, 49, 62, 66, 61, 45, 47, 45, 42, 43, 47, 42, 47, 52, 58, 59, 46, 43, 46, 41, 42, 51, 48, 47, 48, 77, 65, 51, 44, 44, 42, 43, 46, 42, 42, 47, 48, 79, 72, 88, 92, 66, 72, 53, 61, 49, 41, 52, 71, 48, 54, 93, 68, 52, 44, 43, 41, 37, 37, 38, 39, 40, 41, 44, 41, 96, 107, 60, 101, 140, 133, 120, 102, 101, 96, 95, 92, 98, 97, 103, 98, 101, 104, 115, 114, 111, 111, 113, 117, 113, 113, 110, 112, 105, 99, 108, 104, 104, 103, 101, 97, 93, 93, 82, 74, 69, 71, 75, 81, 89, 92, 235, 233, 231, 235, 152, 233, 237, 237, 238, 239, 238, 237, 227, 185, 89, 79, 105, 117, 139, 99, 101, 93, 84, 80, 115, 119, 39, 39, 42, 53, 83, 136, 100, 100, 96, 92, 68, 71, 152, 184, 167, 191, 212, 219, 202, 188, 152, 94, 109, 135, 187, 148, 156, 202, 168, 228, 232, 231, 225, 215, 187, 114, 107, 110, 113, 103, 90, 91, 108, 113, 119, 129, 126, 135, 134, 136, 127, 124, 136, 159, 145, 151, 163, 192, 214, 215, 220, 217, 128, 183, 100, 146, 228, 230, 231, 232, 232, 231, 231, 231, 232, 231, 231, 231, 231, 232, 232, 232, 232, 232, 232, 234, 233, 233, 232, 232, 234, 234, 234, 234, 234, 234, 235, 235, 236, 236, 236, 238, 239, 240, 240, 240, 242, 244, 246, 245, 241, 228, 182, 63, 49, 54, 47, 45, 43, 40, 45, 51, 69, 58, 45, 44, 47, 44, 40, 45, 41, 47, 47, 62, 54, 42, 47, 44, 37, 44, 47, 49, 50, 43, 76, 61, 50, 44, 44, 46, 40, 46, 43, 46, 41, 45, 65, 72, 83, 98, 76, 56, 45, 60, 47, 59, 68, 67, 51, 47, 94, 63, 53, 42, 42, 39, 43, 40, 39, 43, 49, 40, 48, 43, 104, 90, 60, 67, 93, 89, 87, 90, 92, 84, 91, 90, 93, 91, 100, 100, 107, 108, 118, 111, 114, 109, 110, 109, 106, 105, 99, 95, 82, 87, 88, 81, 77, 85, 92, 82, 75, 67, 70, 75, 73, 83, 83, 93, 92, 86, 235, 233, 229, 235, 128, 229, 237, 237, 237, 239, 239, 237, 226, 178, 90, 75, 114, 91, 112, 75, 74, 81, 86, 98, 117, 100, 47, 53, 92, 135, 141, 90, 100, 95, 86, 75, 68, 76, 131, 180, 174, 178, 191, 209, 202, 157, 153, 90, 110, 124, 194, 170, 159, 199, 170, 225, 231, 232, 223, 224, 211, 186, 134, 93, 85, 82, 86, 90, 89, 95, 102, 108, 115, 113, 118, 112, 115, 125, 118, 124, 131, 150, 162, 200, 208, 210, 214, 219, 124, 171, 100, 146, 228, 230, 231, 232, 231, 230, 231, 231, 232, 232, 231, 231, 231, 232, 233, 233, 232, 231, 232, 234, 234, 233, 232, 233, 234, 234, 235, 234, 233, 233, 235, 236, 235, 236, 236, 238, 238, 240, 240, 241, 241, 244, 245, 245, 242, 230, 197, 69, 50, 48, 52, 43, 46, 45, 42, 47, 68, 51, 49, 44, 43, 41, 42, 45, 42, 46, 44, 73, 57, 44, 41, 43, 42, 44, 43, 48, 46, 40, 75, 61, 57, 47, 48, 44, 44, 47, 43, 47, 44, 49, 57, 76, 72, 64, 65, 49, 56, 74, 66, 61, 79, 69, 59, 45, 88, 58, 59, 42, 43, 46, 41, 43, 42, 45, 37, 43, 46, 36, 114, 85, 61, 53, 97, 105, 106, 97, 90, 88, 88, 87, 86, 95, 92, 90, 98, 107, 104, 101, 95, 88, 87, 87, 81, 79, 77, 68, 74, 82, 85, 83, 93, 87, 96, 89, 85, 82, 84, 86, 96, 104, 97, 103, 94, 85, 235, 232, 229, 233, 118, 228, 236, 237, 237, 238, 238, 237, 225, 175, 82, 75, 110, 81, 83, 70, 65, 72, 75, 81, 109, 115, 75, 134, 196, 198, 170, 91, 84, 89, 77, 74, 68, 113, 136, 173, 176, 175, 183, 175, 204, 196, 137, 92, 106, 116, 209, 165, 156, 193, 173, 217, 223, 221, 214, 218, 213, 206, 196, 175, 137, 87, 77, 83, 86, 89, 82, 89, 96, 99, 101, 99, 97, 101, 106, 115, 116, 133, 147, 181, 186, 188, 188, 207, 114, 164, 96, 144, 228, 230, 232, 231, 231, 230, 231, 231, 232, 233, 231, 231, 231, 232, 232, 233, 232, 231, 233, 233, 234, 233, 233, 233, 234, 234, 234, 233, 233, 234, 236, 236, 236, 236, 236, 237, 239, 239, 239, 240, 241, 243, 244, 245, 242, 233, 213, 79, 57, 46, 48, 46, 45, 46, 47, 39, 68, 52, 51, 46, 47, 43, 41, 43, 48, 42, 42, 75, 55, 47, 41, 44, 40, 42, 45, 43, 46, 46, 74, 62, 70, 46, 45, 44, 42, 46, 44, 41, 46, 51, 49, 79, 64, 59, 66, 58, 66, 67, 58, 56, 44, 62, 65, 44, 85, 53, 56, 43, 41, 42, 41, 38, 45, 41, 40, 41, 38, 41, 88, 74, 65, 49, 96, 111, 106, 100, 89, 84, 77, 82, 74, 77, 80, 78, 77, 94, 80, 91, 91, 91, 89, 88, 82, 83, 83, 78, 84, 93, 97, 92, 93, 98, 106, 97, 100, 98, 92, 99, 99, 98, 102, 102, 100, 93, 235, 232, 229, 234, 141, 231, 236, 238, 238, 239, 237, 236, 225, 170, 73, 76, 108, 81, 89, 68, 65, 68, 70, 81, 134, 107, 65, 114, 203, 200, 159, 84, 67, 69, 78, 94, 125, 152, 165, 173, 176, 97, 105, 112, 145, 167, 128, 95, 94, 141, 222, 172, 156, 191, 150, 162, 164, 152, 146, 150, 146, 137, 137, 131, 112, 93, 80, 80, 81, 84, 82, 80, 82, 89, 84, 85, 87, 79, 84, 77, 78, 81, 89, 100, 90, 101, 113, 125, 105, 132, 85, 142, 228, 230, 232, 231, 231, 230, 231, 232, 232, 233, 231, 231, 231, 232, 232, 233, 232, 232, 233, 233, 233, 233, 233, 233, 233, 234, 234, 233, 233, 233, 235, 234, 235, 236, 235, 237, 238, 238, 237, 240, 239, 241, 242, 243, 240, 236, 223, 127, 69, 52, 50, 45, 45, 43, 45, 42, 60, 51, 52, 45, 42, 39, 44, 43, 40, 45, 41, 62, 52, 53, 43, 44, 42, 43, 42, 46, 49, 42, 61, 57, 70, 44, 43, 42, 45, 43, 45, 44, 44, 47, 46, 88, 62, 61, 65, 48, 44, 40, 40, 60, 41, 61, 61, 51, 80, 53, 61, 40, 40, 43, 39, 37, 38, 40, 42, 39, 39, 38, 67, 76, 63, 46, 94, 96, 99, 92, 83, 76, 72, 76, 82, 78, 81, 85, 95, 98, 98, 101, 106, 102, 108, 97, 97, 100, 99, 98, 103, 110, 105, 99, 97, 110, 106, 100, 104, 97, 93, 99, 102, 111, 112, 104, 105, 103, 235, 231, 231, 235, 133, 231, 237, 239, 239, 240, 239, 236, 226, 167, 72, 78, 96, 86, 88, 65, 59, 58, 67, 89, 157, 112, 63, 72, 192, 200, 142, 84, 72, 74, 102, 109, 138, 133, 117, 138, 133, 61, 89, 73, 76, 77, 87, 94, 106, 126, 220, 178, 151, 179, 105, 102, 103, 96, 88, 81, 78, 79, 82, 80, 78, 81, 82, 83, 82, 89, 81, 81, 84, 87, 83, 81, 83, 79, 81, 85, 84, 83, 85, 91, 94, 97, 97, 95, 98, 112, 79, 128, 227, 230, 231, 232, 232, 231, 230, 231, 232, 232, 231, 231, 231, 232, 233, 233, 232, 232, 232, 233, 233, 233, 233, 232, 234, 234, 234, 233, 232, 233, 234, 232, 234, 235, 234, 236, 237, 237, 235, 236, 237, 236, 239, 240, 238, 239, 231, 207, 118, 73, 54, 47, 52, 50, 46, 44, 56, 48, 49, 45, 39, 41, 46, 46, 42, 42, 38, 69, 49, 55, 42, 42, 39, 44, 46, 47, 46, 43, 54, 64, 67, 45, 45, 42, 45, 43, 44, 44, 48, 46, 46, 83, 55, 58, 64, 54, 41, 42, 42, 46, 45, 88, 72, 62, 62, 59, 52, 44, 42, 41, 37, 38, 48, 37, 42, 38, 33, 39, 52, 62, 78, 39, 82, 100, 98, 91, 89, 83, 85, 81, 97, 87, 90, 99, 101, 99, 108, 106, 111, 106, 107, 98, 103, 101, 99, 98, 99, 109, 103, 102, 97, 115, 103, 104, 104, 104, 103, 103, 110, 111, 119, 105, 105, 102, 234, 233, 232, 236, 144, 233, 238, 240, 239, 241, 240, 237, 225, 161, 72, 75, 98, 80, 87, 71, 69, 67, 79, 101, 164, 102, 59, 64, 165, 174, 113, 100, 80, 72, 67, 72, 72, 66, 65, 68, 66, 65, 58, 59, 61, 63, 77, 84, 105, 109, 215, 186, 147, 113, 103, 96, 89, 88, 79, 72, 77, 78, 78, 83, 86, 81, 88, 93, 81, 85, 88, 87, 91, 91, 95, 97, 98, 98, 103, 108, 102, 102, 96, 96, 101, 102, 101, 96, 109, 88, 109, 154, 227, 231, 231, 232, 232, 230, 230, 231, 232, 232, 231, 231, 231, 232, 232, 233, 232, 232, 232, 233, 233, 233, 232, 232, 233, 234, 234, 232, 232, 233, 234, 234, 233, 234, 234, 235, 236, 236, 235, 236, 237, 237, 240, 241, 239, 241, 237, 228, 188, 91, 77, 62, 70, 60, 56, 51, 47, 50, 52, 46, 38, 44, 44, 45, 44, 42, 42, 53, 50, 51, 41, 44, 44, 42, 42, 44, 45, 46, 52, 60, 69, 49, 45, 46, 44, 44, 43, 43, 47, 45, 49, 82, 55, 62, 59, 42, 45, 40, 42, 40, 37, 49, 53, 45, 57, 67, 52, 42, 38, 38, 40, 39, 40, 40, 36, 37, 33, 37, 47, 70, 110, 46, 74, 91, 100, 95, 88, 88, 89, 91, 92, 87, 94, 97, 94, 103, 100, 102, 107, 92, 97, 99, 97, 102, 88, 96, 101, 102, 104, 105, 110, 116, 116, 113, 108, 112, 105, 102, 102, 101, 108, 105, 108, 118, 234, 233, 232, 236, 145, 232, 238, 240, 240, 240, 239, 235, 222, 147, 67, 73, 108, 84, 84, 86, 71, 72, 74, 84, 122, 68, 65, 64, 76, 74, 68, 68, 65, 62, 64, 64, 66, 64, 64, 67, 70, 72, 68, 67, 63, 71, 68, 78, 92, 99, 200, 162, 140, 112, 123, 105, 96, 92, 88, 82, 83, 89, 88, 93, 93, 90, 92, 89, 87, 85, 83, 88, 86, 91, 86, 97, 94, 89, 94, 101, 98, 94, 95, 95, 104, 102, 107, 97, 104, 95, 116, 154, 228, 231, 232, 232, 232, 231, 231, 231, 230, 232, 231, 231, 231, 232, 233, 233, 232, 232, 232, 234, 234, 233, 232, 232, 234, 234, 234, 233, 233, 233, 235, 235, 235, 234, 235, 236, 235, 235, 235, 237, 238, 238, 241, 241, 240, 236, 227, 197, 107, 91, 80, 74, 80, 78, 72, 65, 58, 59, 63, 57, 56, 54, 51, 52, 47, 43, 47, 48, 50, 48, 42, 44, 43, 44, 41, 44, 42, 45, 45, 57, 65, 45, 45, 44, 45, 43, 42, 45, 47, 49, 46, 78, 57, 71, 49, 48, 46, 46, 42, 39, 37, 39, 38, 51, 53, 75, 47, 49, 36, 39, 37, 41, 38, 42, 40, 35, 35, 49, 42, 79, 100, 51, 72, 106, 110, 108, 96, 98, 90, 89, 91, 90, 95, 96, 94, 92, 90, 92, 93, 92, 93, 103, 101, 103, 104, 98, 101, 113, 112, 116, 121, 120, 117, 113, 111, 95, 90, 96, 106, 115, 128, 126, 117, 103, 233, 230, 231, 233, 136, 230, 235, 238, 234, 238, 235, 232, 219, 139, 67, 77, 108, 75, 73, 71, 73, 68, 68, 63, 63, 61, 61, 64, 65, 69, 64, 72, 66, 64, 63, 68, 70, 71, 72, 74, 80, 73, 74, 77, 74, 74, 74, 75, 80, 84, 112, 113, 110, 102, 103, 100, 94, 89, 95, 85, 88, 91, 92, 90, 88, 90, 85, 83, 85, 85, 81, 92, 96, 94, 101, 101, 96, 96, 98, 96, 102, 99, 98, 100, 109, 114, 113, 116, 111, 117, 115, 154, 228, 231, 231, 232, 232, 230, 230, 231, 231, 229, 229, 230, 231, 232, 233, 232, 232, 232, 232, 233, 233, 233, 232, 232, 234, 234, 234, 232, 233, 233, 235, 235, 234, 234, 235, 236, 236, 236, 235, 237, 237, 239, 241, 240, 238, 234, 222, 138, 97, 87, 83, 77, 79, 78, 81, 78, 83, 83, 80, 69, 72, 67, 72, 73, 67, 65, 62, 64, 67, 53, 50, 51, 45, 47, 51, 47, 51, 43, 42, 53, 49, 47, 46, 40, 47, 42, 40, 50, 45, 44, 49, 67, 63, 65, 46, 43, 39, 40, 43, 37, 40, 42, 42, 51, 46, 78, 47, 45, 38, 40, 35, 41, 41, 37, 40, 36, 34, 34, 32, 58, 70, 51, 60, 120, 129, 128, 112, 108, 107, 93, 103, 102, 95, 98, 93, 94, 97, 91, 90, 96, 103, 99, 102, 111, 108, 99, 103, 117, 120, 124, 134, 129, 126, 127, 111, 101, 93, 88, 83, 81, 79, 73, 50, 45, 228, 220, 216, 222, 121, 215, 224, 224, 221, 221, 221, 213, 201, 119, 73, 72, 85, 67, 69, 69, 67, 65, 70, 72, 63, 67, 65, 71, 73, 70, 68, 70, 70, 72, 71, 74, 75, 70, 69, 76, 71, 72, 70, 82, 80, 86, 86, 90, 102, 109, 180, 185, 134, 111, 107, 107, 114, 106, 103, 99, 99, 97, 96, 100, 102, 93, 89, 93, 97, 94, 94, 98, 101, 93, 103, 92, 95, 96, 99, 100, 103, 102, 107, 105, 111, 122, 122, 138, 114, 130, 119, 152, 229, 231, 231, 232, 232, 231, 231, 231, 232, 231, 232, 230, 231, 231, 233, 233, 231, 232, 232, 233, 233, 232, 232, 232, 233, 234, 233, 233, 233, 233, 234, 235, 235, 233, 235, 236, 237, 236, 236, 237, 236, 240, 242, 239, 236, 229, 208, 107, 95, 84, 82, 78, 82, 79, 74, 75, 93, 84, 78, 75, 77, 72, 70, 67, 71, 72, 75, 69, 76, 69, 73, 66, 69, 68, 67, 66, 62, 61, 57, 59, 62, 54, 50, 48, 49, 47, 56, 44, 49, 53, 48, 56, 75, 71, 49, 44, 43, 40, 39, 41, 41, 36, 44, 45, 43, 71, 49, 48, 38, 39, 39, 46, 36, 38, 38, 36, 32, 33, 37, 51, 52, 57, 50, 108, 116, 110, 107, 106, 101, 97, 103, 103, 93, 101, 93, 101, 103, 104, 107, 108, 116, 121, 124, 121, 129, 115, 114, 114, 114, 102, 88, 83, 77, 65, 58, 50, 46, 44, 48, 49, 39, 63, 37, 36, 204, 200, 200, 202, 114, 200, 206, 197, 204, 204, 204, 201, 195, 114, 68, 69, 72, 67, 64, 66, 67, 73, 67, 68, 70, 79, 71, 76, 69, 67, 69, 74, 73, 68, 72, 71, 78, 77, 76, 81, 86, 91, 87, 88, 88, 86, 90, 89, 107, 109, 190, 200, 137, 122, 108, 113, 114, 112, 107, 112, 106, 110, 105, 103, 107, 96, 97, 99, 97, 99, 106, 93, 98, 102, 105, 99, 100, 104, 108, 105, 105, 108, 108, 118, 126, 132, 157, 181, 118, 143, 117, 160, 229, 230, 231, 232, 231, 231, 231, 231, 232, 232, 231, 231, 231, 232, 232, 232, 231, 232, 232, 233, 233, 232, 232, 232, 233, 234, 234, 233, 233, 233, 234, 235, 235, 234, 235, 236, 237, 236, 236, 237, 237, 240, 240, 240, 236, 227, 200, 106, 89, 86, 79, 80, 81, 83, 82, 76, 96, 88, 89, 76, 73, 71, 75, 77, 71, 71, 74, 78, 85, 78, 69, 74, 69, 74, 73, 75, 74, 73, 77, 70, 75, 76, 65, 65, 58, 69, 66, 62, 62, 63, 67, 81, 100, 96, 69, 57, 54, 46, 40, 47, 44, 41, 43, 45, 41, 62, 49, 52, 39, 39, 43, 37, 37, 40, 39, 37, 37, 37, 49, 48, 61, 54, 44, 98, 126, 120, 115, 108, 111, 103, 107, 109, 96, 104, 105, 109, 107, 105, 103, 95, 100, 95, 87, 85, 74, 66, 59, 58, 61, 50, 44, 44, 43, 39, 40, 36, 38, 37, 38, 50, 45, 45, 44, 54, 207, 209, 205, 208, 105, 207, 208, 214, 212, 210, 211, 207, 201, 108, 72, 73, 73, 69, 68, 68, 68, 68, 65, 66, 67, 69, 74, 74, 72, 79, 78, 74, 79, 71, 80, 77, 80, 81, 82, 89, 88, 89, 82, 93, 94, 92, 88, 93, 104, 123, 188, 179, 140, 173, 128, 140, 142, 141, 137, 141, 137, 138, 133, 129, 114, 100, 102, 100, 102, 100, 102, 103, 112, 104, 105, 110, 112, 116, 113, 122, 122, 130, 137, 163, 170, 178, 196, 209, 134, 158, 125, 156, 229, 231, 232, 231, 231, 231, 230, 231, 231, 232, 230, 231, 232, 232, 233, 233, 231, 232, 232, 233, 233, 233, 232, 232, 233, 234, 233, 232, 233, 233, 234, 235, 234, 234, 234, 236, 236, 236, 235, 235, 237, 240, 238, 238, 235, 225, 192, 98, 98, 89, 81, 81, 83, 86, 84, 76, 105, 86, 85, 76, 75, 74, 75, 72, 78, 79, 78, 85, 93, 80, 74, 75, 76, 71, 72, 75, 74, 78, 69, 84, 76, 77, 73, 73, 68, 78, 78, 73, 72, 68, 75, 79, 91, 73, 64, 64, 62, 55, 51, 52, 56, 48, 56, 51, 44, 53, 48, 50, 42, 39, 37, 36, 39, 42, 45, 40, 41, 43, 42, 48, 57, 53, 55, 73, 108, 95, 86, 65, 68, 71, 67, 72, 70, 64, 58, 59, 58, 50, 53, 50, 46, 50, 47, 43, 50, 41, 43, 45, 40, 43, 49, 48, 47, 48, 50, 44, 50, 49, 54, 54, 55, 56, 54, 55, 205, 208, 208, 208, 121, 208, 211, 215, 214, 213, 210, 210, 199, 134, 80, 67, 69, 76, 72, 71, 68, 71, 73, 71, 73, 76, 75, 76, 83, 82, 81, 78, 78, 75, 82, 86, 84, 83, 90, 92, 96, 94, 98, 104, 107, 114, 106, 92, 107, 124, 195, 171, 146, 190, 156, 180, 181, 175, 177, 181, 177, 169, 160, 138, 114, 100, 103, 103, 105, 109, 109, 114, 119, 117, 120, 123, 117, 119, 125, 128, 131, 145, 146, 168, 180, 185, 209, 212, 132, 159, 127, 162, 229, 230, 232, 231, 231, 231, 230, 231, 232, 232, 231, 231, 231, 232, 232, 233, 231, 232, 232, 233, 233, 233, 232, 232, 234, 233, 233, 233, 233, 233, 233, 234, 233, 233, 233, 235, 236, 236, 234, 235, 236, 239, 238, 237, 234, 224, 184, 96, 91, 90, 91, 87, 85, 86, 83, 84, 104, 85, 85, 76, 76, 82, 78, 81, 83, 87, 77, 91, 92, 82, 77, 74, 73, 78, 79, 76, 80, 74, 84, 90, 89, 83, 79, 78, 73, 80, 70, 77, 71, 72, 70, 81, 101, 100, 80, 74, 74, 69, 73, 68, 67, 64, 68, 69, 62, 55, 55, 50, 46, 44, 44, 37, 45, 44, 45, 47, 43, 46, 55, 65, 75, 88, 107, 88, 75, 57, 59, 42, 42, 44, 44, 51, 46, 41, 41, 42, 40, 42, 43, 45, 41, 43, 47, 47, 48, 52, 51, 59, 70, 70, 77, 72, 74, 74, 67, 62, 64, 66, 68, 66, 72, 62, 60, 60, 199, 206, 205, 209, 120, 206, 209, 212, 213, 210, 208, 207, 197, 115, 87, 84, 82, 83, 83, 74, 77, 78, 81, 85, 83, 87, 83, 84, 94, 96, 84, 84, 78, 82, 82, 91, 99, 102, 112, 132, 126, 99, 117, 129, 151, 152, 127, 103, 121, 123, 173, 201, 156, 197, 160, 185, 189, 187, 188, 181, 175, 145, 127, 116, 110, 109, 112, 107, 107, 115, 117, 114, 126, 129, 128, 129, 129, 130, 135, 146, 143, 145, 148, 172, 180, 188, 211, 209, 128, 158, 121, 160, 229, 231, 232, 232, 231, 230, 231, 231, 231, 232, 231, 231, 232, 232, 232, 233, 232, 231, 232, 233, 233, 233, 232, 232, 234, 234, 233, 233, 233, 233, 233, 234, 233, 233, 234, 234, 236, 237, 233, 235, 236, 239, 237, 236, 233, 224, 179, 104, 94, 96, 87, 86, 84, 82, 84, 81, 111, 87, 87, 81, 78, 80, 71, 81, 84, 80, 80, 92, 88, 88, 83, 79, 79, 76, 79, 81, 77, 84, 76, 91, 88, 83, 75, 75, 72, 75, 79, 80, 74, 71, 81, 78, 102, 88, 80, 75, 72, 70, 74, 66, 69, 77, 76, 76, 68, 70, 68, 69, 66, 63, 61, 53, 58, 55, 58, 54, 53, 51, 70, 88, 117, 134, 132, 139, 93, 73, 60, 41, 46, 44, 50, 44, 51, 52, 56, 58, 50, 55, 53, 55, 59, 66, 67, 57, 63, 60, 64, 75, 72, 74, 80, 85, 86, 90, 83, 77, 80, 81, 83, 94, 98, 99, 99, 102, 202, 204, 204, 210, 130, 207, 209, 210, 214, 212, 208, 203, 195, 113, 85, 88, 83, 91, 90, 84, 85, 87, 79, 83, 96, 81, 90, 94, 121, 121, 104, 98, 92, 89, 99, 110, 120, 130, 137, 148, 142, 140, 147, 156, 169, 144, 129, 96, 122, 132, 158, 195, 159, 188, 157, 189, 191, 191, 184, 176, 147, 116, 122, 126, 123, 119, 116, 116, 121, 123, 127, 129, 130, 130, 135, 136, 129, 132, 138, 149, 147, 149, 154, 170, 181, 186, 208, 202, 126, 159, 123, 158, 228, 229, 231, 232, 231, 231, 230, 231, 232, 232, 231, 231, 231, 232, 232, 232, 232, 231, 232, 233, 233, 232, 232, 232, 233, 234, 233, 232, 233, 233, 233, 234, 234, 232, 234, 235, 237, 236, 234, 236, 237, 238, 236, 235, 233, 224, 172, 103, 100, 94, 97, 87, 91, 91, 90, 91, 107, 87, 84, 77, 74, 79, 71, 76, 80, 81, 76, 96, 89, 83, 79, 77, 80, 73, 76, 77, 70, 76, 79, 96, 95, 83, 77, 77, 74, 75, 81, 76, 79, 76, 79, 81, 97, 90, 79, 78, 73, 75, 71, 70, 71, 73, 71, 68, 70, 86, 86, 71, 74, 65, 64, 73, 69, 64, 64, 68, 63, 65, 66, 80, 110, 112, 103, 129, 107, 97, 83, 49, 53, 56, 60, 58, 64, 59, 61, 68, 66, 64, 76, 70, 74, 84, 83, 82, 89, 92, 92, 92, 106, 104, 104, 100, 108, 102, 96, 99, 97, 97, 98, 100, 103, 107, 100, 100, 201, 201, 200, 205, 129, 200, 208, 209, 211, 208, 203, 199, 195, 108, 95, 93, 97, 88, 90, 89, 108, 87, 96, 97, 137, 89, 86, 96, 152, 151, 108, 90, 88, 100, 93, 100, 107, 122, 135, 149, 143, 151, 160, 176, 160, 136, 126, 97, 117, 132, 151, 173, 155, 190, 160, 191, 187, 177, 173, 152, 122, 128, 137, 131, 121, 125, 123, 123, 132, 135, 132, 136, 136, 134, 143, 140, 135, 136, 145, 144, 153, 157, 153, 169, 184, 188, 212, 195, 125, 160, 127, 155, 227, 229, 231, 232, 231, 231, 230, 231, 231, 232, 231, 231, 232, 232, 233, 233, 232, 231, 232, 233, 233, 232, 232, 232, 233, 234, 233, 232, 233, 232, 234, 234, 233, 233, 233, 235, 236, 235, 233, 234, 235, 237, 236, 235, 231, 221, 166, 108, 102, 96, 98, 90, 91, 91, 90, 92, 118, 98, 82, 85, 82, 83, 75, 83, 80, 83, 80, 96, 86, 85, 81, 78, 79, 75, 79, 80, 85, 76, 81, 103, 100, 83, 81, 77, 75, 81, 78, 80, 75, 77, 81, 85, 98, 91, 85, 77, 76, 72, 81, 75, 74, 73, 69, 74, 68, 93, 84, 74, 73, 65, 68, 69, 65, 64, 70, 70, 64, 69, 76, 84, 104, 109, 104, 116, 103, 94, 83, 62, 60, 64, 70, 65, 73, 74, 79, 92, 95, 101, 112, 110, 115, 115, 109, 110, 104, 106, 103, 100, 105, 108, 106, 102, 104, 104, 95, 100, 100, 103, 103, 105, 105, 104, 99, 102, 204, 200, 203, 206, 140, 202, 210, 211, 210, 204, 204, 200, 188, 108, 94, 101, 95, 97, 98, 97, 94, 97, 95, 105, 149, 88, 88, 112, 165, 160, 111, 97, 94, 96, 97, 91, 94, 112, 136, 156, 139, 154, 171, 175, 167, 155, 126, 99, 128, 149, 169, 161, 166, 191, 161, 184, 184, 149, 156, 131, 127, 128, 131, 135, 135, 146, 137, 138, 139, 141, 137, 143, 139, 141, 145, 138, 138, 143, 146, 145, 148, 156, 160, 168, 191, 193, 215, 188, 126, 158, 124, 152, 227, 231, 231, 231, 232, 231, 230, 231, 232, 232, 231, 231, 231, 232, 233, 233, 232, 232, 231, 233, 233, 232, 232, 232, 233, 234, 233, 233, 232, 231, 234, 234, 233, 234, 234, 236, 236, 235, 233, 234, 233, 236, 236, 232, 231, 221, 157, 103, 106, 95, 94, 92, 91, 92, 89, 93, 115, 95, 91, 86, 78, 81, 86, 84, 80, 81, 77, 99, 89, 83, 84, 82, 82, 79, 82, 79, 81, 76, 88, 99, 97, 82, 76, 82, 80, 82, 80, 76, 81, 74, 80, 94, 97, 93, 84, 79, 78, 78, 79, 75, 78, 71, 75, 76, 80, 99, 90, 82, 70, 76, 65, 72, 68, 62, 69, 72, 69, 74, 75, 80, 89, 99, 112, 103, 94, 91, 79, 79, 73, 79, 97, 101, 105, 102, 111, 106, 102, 109, 107, 107, 107, 109, 109, 101, 103, 106, 111, 107, 105, 102, 103, 107, 109, 101, 98, 100, 99, 98, 98, 100, 102, 101, 98, 100, 202, 203, 202, 205, 129, 205, 208, 209, 205, 206, 204, 196, 191, 112, 94, 96, 97, 94, 100, 92, 92, 96, 96, 101, 142, 88, 94, 132, 164, 160, 116, 103, 102, 101, 96, 97, 103, 103, 144, 153, 147, 173, 181, 179, 176, 158, 139, 100, 131, 154, 170, 153, 161, 187, 165, 179, 179, 151, 146, 134, 141, 143, 148, 150, 155, 149, 141, 140, 147, 143, 139, 145, 140, 144, 143, 142, 139, 140, 139, 146, 153, 153, 158, 171, 189, 191, 208, 176, 130, 159, 124, 153, 226, 230, 230, 232, 231, 230, 230, 231, 231, 232, 231, 231, 231, 232, 232, 232, 232, 232, 232, 233, 233, 232, 232, 232, 233, 234, 233, 232, 232, 232, 234, 233, 233, 234, 234, 234, 235, 233, 231, 234, 234, 237, 237, 231, 231, 219, 149, 109, 103, 97, 98, 101, 96, 90, 93, 97, 108, 96, 89, 84, 81, 84, 86, 85, 85, 80, 81, 96, 82, 84, 85, 84, 90, 85, 82, 82, 90, 83, 92, 98, 98, 89, 80, 80, 83, 83, 81, 80, 77, 77, 86, 99, 104, 94, 90, 97, 78, 79, 83, 76, 80, 82, 87, 85, 82, 93, 87, 87, 78, 76, 69, 77, 69, 75, 73, 72, 74, 67, 84, 72, 90, 84, 95, 93, 109, 110, 103, 98, 102, 107, 107, 107, 101, 107, 105, 100, 104, 102, 99, 100, 102, 109, 105, 103, 98, 99, 106, 105, 105, 103, 102, 103, 107, 107, 106, 101, 107, 103, 103, 97, 101, 108, 103, 103, 201, 202, 200, 204, 138, 206, 212, 210, 205, 205, 208, 200, 191, 106, 97, 94, 94, 98, 102, 97, 96, 98, 96, 102, 137, 94, 95, 135, 153, 153, 111, 106, 109, 107, 100, 100, 100, 110, 162, 160, 151, 174, 183, 180, 175, 162, 139, 103, 129, 150, 163, 152, 156, 188, 161, 182, 176, 155, 153, 147, 149, 155, 157, 163, 161, 150, 144, 145, 147, 143, 142, 146, 144, 146, 146, 145, 145, 145, 142, 154, 158, 164, 165, 176, 190, 194, 199, 158, 125, 155, 126, 154, 227, 230, 231, 231, 231, 230, 230, 230, 232, 232, 231, 231, 231, 232, 232, 232, 232, 232, 232, 233, 233, 233, 232, 231, 233, 234, 233, 232, 230, 232, 234, 231, 233, 232, 233, 232, 235, 231, 231, 231, 232, 232, 236, 229, 227, 218, 148, 116, 113, 114, 104, 109, 104, 101, 101, 103, 116, 103, 88, 88, 83, 82, 83, 84, 79, 87, 85, 99, 94, 86, 86, 87, 89, 91, 84, 89, 86, 86, 90, 102, 95, 87, 81, 83, 84, 85, 82, 82, 90, 85, 88, 105, 107, 95, 100, 93, 92, 87, 84, 81, 83, 79, 96, 99, 94, 112, 91, 94, 83, 81, 78, 79, 79, 78, 81, 75, 81, 80, 80, 78, 98, 89, 88, 90, 107, 114, 109, 105, 114, 106, 106, 105, 107, 104, 101, 110, 102, 109, 99, 105, 102, 102, 107, 102, 99, 102, 104, 106, 101, 104, 104, 99, 105, 103, 101, 99, 106, 106, 96, 101, 101, 102, 100, 105, 199, 204, 203, 204, 146, 203, 210, 208, 208, 203, 203, 197, 186, 113, 96, 94, 94, 95, 104, 99, 97, 99, 93, 103, 127, 94, 83, 93, 103, 109, 115, 109, 109, 115, 111, 102, 109, 134, 168, 164, 164, 172, 177, 182, 172, 167, 137, 100, 130, 156, 162, 149, 160, 184, 164, 184, 184, 155, 156, 155, 165, 165, 167, 171, 169, 151, 144, 148, 150, 146, 148, 142, 147, 144, 140, 152, 152, 162, 155, 158, 156, 157, 167, 176, 192, 195, 191, 154, 129, 157, 125, 152, 227, 230, 231, 231, 231, 231, 230, 231, 232, 232, 232, 231, 231, 232, 233, 233, 232, 231, 232, 233, 233, 233, 232, 231, 232, 231, 232, 232, 227, 229, 231, 230, 231, 231, 231, 232, 234, 232, 232, 229, 228, 231, 234, 231, 225, 219, 151, 113, 113, 114, 107, 109, 110, 101, 106, 105, 116, 102, 99, 91, 91, 90, 88, 92, 85, 88, 90, 97, 96, 99, 86, 89, 90, 92, 85, 88, 86, 92, 92, 106, 102, 95, 81, 82, 89, 84, 86, 84, 87, 85, 96, 103, 99, 108, 97, 98, 92, 90, 91, 84, 91, 85, 105, 106, 92, 109, 89, 95, 87, 89, 80, 84, 83, 85, 89, 91, 84, 83, 83, 86, 115, 97, 97, 100, 113, 118, 111, 109, 106, 109, 106, 111, 108, 115, 109, 106, 105, 113, 102, 111, 106, 113, 114, 110, 106, 106, 105, 104, 109, 105, 99, 101, 103, 103, 96, 99, 99, 98, 94, 101, 102, 96, 101, 99, 197, 201, 199, 203, 132, 198, 206, 207, 208, 204, 200, 196, 182, 104, 104, 100, 91, 102, 107, 103, 99, 104, 106, 104, 124, 87, 84, 77, 87, 81, 126, 122, 115, 107, 105, 96, 105, 141, 164, 161, 159, 170, 180, 180, 171, 167, 137, 102, 131, 153, 159, 140, 162, 179, 171, 185, 182, 159, 152, 159, 169, 164, 165, 167, 163, 148, 144, 144, 141, 140, 140, 142, 136, 140, 139, 144, 153, 161, 159, 166, 164, 167, 168, 175, 194, 190, 177, 149, 139, 155, 132, 160, 228, 230, 231, 231, 231, 230, 230, 231, 232, 232, 231, 231, 231, 232, 233, 232, 232, 231, 232, 233, 233, 232, 231, 231, 232, 231, 232, 231, 226, 229, 231, 230, 229, 232, 230, 231, 231, 233, 232, 228, 227, 232, 233, 228, 227, 216, 150, 117, 119, 122, 113, 115, 115, 109, 110, 110, 116, 107, 98, 92, 98, 86, 93, 95, 94, 97, 92, 103, 100, 94, 96, 86, 90, 93, 87, 85, 87, 84, 97, 99, 104, 98, 87, 88, 93, 86, 90, 89, 90, 95, 94, 105, 96, 105, 100, 103, 95, 100, 93, 89, 97, 97, 98, 104, 89, 112, 96, 99, 89, 85, 86, 82, 87, 87, 85, 87, 85, 83, 87, 95, 108, 109, 94, 100, 113, 117, 114, 108, 108, 104, 108, 107, 110, 117, 110, 115, 108, 107, 108, 104, 109, 109, 111, 104, 102, 106, 100, 101, 107, 104, 110, 103, 100, 107, 101, 103, 93, 101, 99, 101, 97, 94, 94, 95, 198, 199, 197, 200, 144, 195, 208, 206, 210, 208, 197, 197, 180, 107, 104, 102, 93, 109, 108, 96, 101, 99, 100, 110, 125, 95, 83, 80, 90, 85, 119, 137, 124, 111, 106, 112, 124, 142, 175, 157, 162, 168, 174, 178, 171, 165, 139, 106, 138, 145, 153, 136, 164, 181, 178, 183, 182, 166, 152, 145, 148, 143, 144, 140, 137, 134, 130, 129, 131, 129, 122, 131, 122, 128, 140, 144, 147, 152, 161, 163, 163, 167, 169, 178, 191, 193, 171, 148, 139, 161, 133, 158, 228, 230, 232, 232, 231, 231, 231, 231, 232, 232, 231, 231, 230, 232, 232, 232, 232, 231, 231, 232, 233, 233, 231, 231, 231, 232, 232, 231, 228, 230, 232, 229, 226, 231, 230, 231, 233, 232, 229, 230, 227, 231, 234, 229, 223, 215, 144, 124, 142, 125, 124, 120, 119, 113, 112, 112, 117, 107, 100, 103, 100, 95, 92, 95, 98, 103, 96, 104, 101, 89, 96, 91, 93, 90, 86, 91, 96, 86, 104, 103, 105, 94, 95, 86, 91, 89, 91, 89, 86, 92, 97, 112, 100, 110, 109, 95, 94, 99, 104, 101, 97, 97, 107, 102, 102, 109, 102, 97, 91, 92, 86, 84, 88, 93, 91, 93, 82, 87, 88, 97, 110, 113, 89, 102, 111, 109, 108, 102, 108, 101, 109, 112, 112, 114, 110, 113, 114, 111, 104, 105, 103, 110, 113, 107, 106, 103, 103, 103, 110, 105, 106, 107, 102, 101, 102, 102, 104, 105, 103, 103, 105, 98, 107, 106, 201, 196, 197, 203, 127, 200, 207, 208, 205, 208, 203, 191, 175, 107, 102, 108, 99, 115, 110, 100, 101, 102, 104, 115, 125, 96, 85, 85, 86, 88, 116, 134, 137, 125, 120, 126, 138, 156, 155, 151, 156, 159, 176, 175, 169, 168, 145, 106, 128, 144, 166, 141, 156, 184, 172, 178, 179, 178, 161, 150, 144, 138, 138, 137, 133, 130, 126, 124, 126, 123, 126, 123, 131, 133, 136, 142, 148, 156, 160, 162, 170, 167, 172, 180, 191, 189, 169, 155, 141, 156, 135, 166, 228, 230, 232, 232, 231, 230, 230, 230, 232, 232, 231, 231, 230, 232, 232, 232, 231, 231, 232, 232, 233, 232, 231, 231, 231, 231, 231, 230, 228, 229, 230, 228, 228, 230, 229, 231, 230, 230, 228, 228, 227, 229, 229, 227, 220, 216, 144, 127, 144, 125, 121, 119, 118, 117, 115, 115, 119, 114, 107, 103, 100, 101, 97, 101, 99, 104, 103, 105, 102, 97, 95, 93, 89, 93, 94, 96, 89, 96, 102, 108, 105, 101, 94, 97, 91, 95, 90, 92, 93, 89, 94, 110, 105, 108, 102, 102, 103, 93, 107, 106, 100, 108, 109, 101, 97, 118, 101, 98, 103, 91, 87, 91, 90, 91, 94, 93, 91, 90, 98, 101, 117, 120, 95, 106, 108, 115, 114, 104, 104, 113, 111, 115, 110, 110, 109, 108, 114, 112, 108, 112, 110, 115, 110, 117, 111, 108, 113, 102, 113, 113, 102, 110, 112, 110, 109, 108, 107, 110, 107, 109, 110, 103, 115, 110, 196, 198, 200, 204, 118, 202, 207, 205, 211, 205, 201, 191, 174, 109, 102, 102, 100, 122, 106, 104, 102, 114, 109, 123, 125, 102, 87, 82, 84, 93, 118, 134, 128, 111, 110, 115, 110, 130, 120, 130, 133, 140, 172, 175, 168, 172, 141, 105, 134, 148, 179, 148, 156, 167, 169, 184, 181, 184, 172, 166, 157, 157, 157, 154, 149, 142, 134, 136, 134, 128, 128, 131, 132, 135, 143, 144, 159, 162, 172, 171, 170, 173, 175, 186, 193, 189, 167, 154, 140, 153, 140, 169, 228, 230, 232, 232, 231, 231, 230, 230, 232, 231, 231, 231, 231, 232, 232, 232, 231, 231, 231, 232, 232, 231, 231, 230, 231, 230, 229, 229, 227, 228, 229, 228, 228, 225, 225, 230, 229, 230, 227, 227, 226, 227, 228, 227, 219, 214, 150, 126, 131, 128, 127, 121, 120, 121, 120, 118, 120, 116, 114, 112, 105, 103, 102, 104, 105, 107, 106, 112, 105, 100, 94, 93, 98, 93, 96, 94, 100, 95, 100, 110, 104, 98, 98, 99, 99, 97, 95, 98, 94, 97, 108, 118, 104, 108, 113, 99, 103, 97, 94, 94, 100, 110, 103, 107, 99, 113, 101, 100, 90, 90, 87, 90, 91, 89, 95, 94, 92, 92, 96, 112, 122, 124, 101, 110, 120, 123, 119, 107, 104, 110, 102, 113, 114, 116, 115, 117, 118, 117, 123, 122, 120, 117, 124, 117, 116, 119, 112, 108, 116, 116, 110, 112, 111, 112, 106, 111, 104, 108, 111, 110, 111, 105, 113, 112, 202, 202, 200, 203, 139, 205, 208, 205, 207, 203, 203, 196, 176, 111, 100, 106, 98, 116, 112, 110, 107, 111, 114, 120, 125, 114, 92, 85, 89, 89, 117, 135, 121, 106, 109, 106, 101, 108, 116, 132, 136, 128, 166, 167, 172, 169, 138, 112, 133, 154, 177, 138, 161, 155, 173, 190, 187, 190, 187, 177, 179, 169, 171, 171, 161, 159, 147, 149, 141, 135, 134, 137, 151, 148, 140, 155, 160, 171, 176, 176, 178, 181, 179, 192, 191, 189, 172, 144, 141, 157, 139, 168, 228, 230, 232, 232, 231, 230, 230, 231, 232, 231, 231, 231, 231, 232, 232, 232, 231, 231, 231, 232, 232, 231, 230, 228, 229, 227, 230, 228, 228, 228, 230, 228, 228, 227, 224, 226, 229, 231, 228, 228, 226, 226, 227, 223, 219, 213, 151, 130, 126, 131, 127, 124, 130, 125, 115, 128, 127, 118, 115, 110, 107, 100, 102, 103, 110, 106, 107, 117, 108, 100, 99, 98, 101, 103, 93, 92, 96, 96, 100, 105, 107, 102, 97, 98, 95, 100, 97, 97, 98, 97, 100, 120, 107, 111, 111, 108, 107, 97, 117, 104, 102, 104, 116, 102, 100, 126, 105, 104, 96, 95, 96, 95, 96, 98, 95, 92, 98, 95, 101, 113, 124, 125, 98, 115, 118, 118, 115, 107, 111, 111, 117, 112, 119, 114, 118, 112, 118, 118, 127, 120, 120, 116, 120, 117, 120, 119, 112, 110, 114, 109, 113, 119, 114, 113, 115, 105, 107, 108, 112, 105, 110, 113, 111, 114, 200, 201, 201, 199, 128, 204, 205, 203, 204, 199, 202, 196, 165, 110, 94, 108, 104, 113, 112, 117, 114, 114, 123, 119, 129, 117, 96, 88, 91, 91, 120, 131, 111, 114, 118, 108, 102, 105, 111, 129, 130, 124, 140, 165, 166, 165, 138, 116, 140, 148, 178, 138, 151, 151, 174, 191, 189, 191, 189, 188, 189, 183, 184, 183, 174, 172, 164, 160, 154, 139, 137, 138, 159, 162, 170, 180, 177, 182, 189, 191, 193, 196, 196, 202, 192, 190, 167, 147, 137, 152, 135, 163, 227, 230, 231, 232, 232, 230, 230, 231, 232, 232, 232, 231, 231, 232, 232, 231, 231, 231, 230, 231, 232, 228, 230, 227, 228, 228, 230, 228, 227, 229, 228, 227, 227, 225, 225, 228, 228, 230, 223, 226, 226, 220, 226, 223, 219, 213, 146, 134, 132, 131, 133, 123, 125, 123, 121, 124, 128, 119, 115, 114, 113, 106, 106, 105, 105, 105, 103, 113, 113, 105, 105, 99, 101, 105, 101, 95, 99, 105, 104, 110, 109, 105, 106, 98, 101, 107, 101, 102, 103, 105, 103, 120, 110, 111, 117, 100, 103, 100, 119, 104, 108, 106, 116, 107, 103, 123, 107, 103, 101, 98, 103, 97, 94, 100, 99, 102, 91, 96, 104, 116, 124, 115, 103, 116, 118, 121, 122, 115, 114, 112, 115, 116, 115, 111, 114, 112, 118, 117, 113, 116, 116, 118, 124, 121, 114, 116, 115, 110, 114, 109, 112, 110, 114, 116, 116, 111, 107, 113, 112, 110, 111, 111, 115, 109, 198, 198, 196, 203, 126, 200, 202, 204, 201, 202, 198, 197, 159, 114, 106, 112, 110, 122, 115, 121, 113, 111, 118, 122, 133, 129, 108, 97, 98, 103, 120, 131, 130, 130, 132, 117, 113, 109, 119, 129, 139, 118, 123, 147, 157, 161, 138, 121, 135, 150, 176, 134, 151, 148, 174, 188, 185, 189, 191, 190, 187, 187, 190, 188, 187, 181, 177, 165, 157, 147, 144, 140, 160, 172, 183, 190, 196, 196, 198, 204, 201, 204, 203, 206, 198, 192, 163, 150, 142, 147, 136, 162, 226, 230, 231, 232, 231, 230, 230, 231, 232, 231, 232, 230, 231, 231, 231, 231, 230, 231, 231, 231, 229, 226, 228, 229, 228, 228, 230, 227, 225, 225, 226, 228, 225, 223, 225, 224, 224, 228, 225, 227, 225, 224, 225, 224, 219, 213, 148, 138, 132, 130, 127, 130, 129, 126, 126, 130, 125, 122, 114, 114, 115, 112, 110, 110, 116, 110, 107, 115, 113, 112, 109, 106, 108, 106, 106, 103, 99, 105, 105, 111, 108, 111, 109, 104, 108, 103, 103, 107, 105, 106, 103, 122, 105, 114, 114, 109, 111, 108, 118, 110, 116, 111, 118, 117, 105, 130, 112, 108, 105, 101, 105, 102, 98, 100, 99, 99, 98, 101, 108, 121, 121, 125, 103, 112, 122, 116, 111, 116, 112, 116, 115, 117, 112, 120, 122, 118, 120, 121, 124, 120, 125, 126, 124, 120, 122, 115, 115, 115, 119, 117, 115, 106, 115, 111, 113, 111, 109, 120, 113, 111, 116, 112, 113, 113, 197, 193, 193, 199, 124, 199, 202, 201, 202, 198, 199, 192, 155, 108, 105, 109, 117, 131, 116, 115, 122, 117, 124, 135, 145, 141, 112, 102, 102, 112, 121, 142, 158, 156, 154, 129, 128, 123, 123, 121, 122, 121, 120, 124, 154, 158, 140, 121, 135, 148, 168, 142, 149, 148, 173, 186, 189, 189, 189, 191, 190, 190, 194, 192, 189, 190, 187, 176, 160, 152, 146, 145, 152, 179, 192, 194, 196, 203, 198, 209, 207, 207, 205, 206, 197, 189, 161, 154, 143, 153, 133, 161, 224, 230, 231, 230, 230, 229, 230, 230, 231, 231, 231, 231, 231, 231, 232, 232, 231, 231, 231, 231, 231, 226, 228, 225, 228, 228, 230, 226, 226, 226, 227, 228, 226, 223, 224, 224, 225, 225, 225, 225, 223, 225, 225, 223, 220, 217, 152, 138, 134, 129, 129, 126, 131, 126, 125, 126, 131, 122, 114, 114, 112, 106, 111, 112, 113, 112, 107, 118, 115, 110, 109, 108, 110, 104, 104, 114, 105, 109, 107, 113, 115, 112, 107, 104, 110, 109, 107, 112, 107, 106, 106, 127, 116, 115, 117, 115, 115, 111, 115, 107, 115, 107, 122, 112, 106, 132, 110, 113, 103, 102, 102, 107, 101, 104, 112, 106, 102, 101, 106, 123, 120, 119, 103, 119, 113, 118, 120, 120, 112, 120, 123, 121, 117, 121, 118, 122, 124, 123, 124, 118, 120, 122, 123, 116, 125, 119, 112, 118, 116, 115, 118, 111, 113, 114, 115, 112, 108, 109, 111, 118, 115, 114, 114, 115, 198, 192, 191, 194, 135, 198, 198, 198, 202, 197, 195, 190, 151, 111, 109, 117, 122, 137, 122, 120, 134, 124, 131, 133, 156, 146, 105, 101, 104, 124, 125, 152, 165, 165, 158, 135, 127, 125, 128, 118, 109, 113, 113, 123, 139, 158, 141, 111, 132, 150, 153, 136, 149, 144, 175, 192, 192, 195, 193, 190, 191, 194, 195, 192, 193, 193, 192, 185, 176, 152, 150, 150, 149, 180, 191, 192, 198, 201, 201, 206, 204, 205, 204, 203, 191, 190, 164, 161, 142, 156, 144, 162, 223, 230, 231, 231, 231, 230, 230, 231, 232, 230, 230, 230, 231, 232, 231, 230, 230, 230, 230, 231, 230, 229, 228, 224, 227, 230, 230, 227, 227, 227, 229, 224, 224, 224, 222, 225, 224, 225, 225, 226, 226, 224, 223, 223, 221, 212, 162, 137, 135, 129, 133, 127, 132, 129, 126, 126, 129, 125, 125, 113, 115, 110, 109, 117, 112, 105, 109, 120, 113, 114, 113, 106, 108, 113, 106, 102, 105, 108, 106, 116, 115, 110, 106, 108, 112, 109, 111, 103, 105, 108, 106, 124, 112, 117, 115, 115, 117, 117, 115, 114, 114, 115, 121, 117, 112, 134, 117, 117, 110, 119, 115, 101, 104, 107, 110, 105, 125, 109, 111, 125, 120, 123, 108, 122, 117, 118, 123, 115, 121, 118, 117, 123, 123, 114, 125, 125, 125, 124, 121, 122, 125, 126, 122, 123, 124, 120, 117, 120, 113, 114, 122, 108, 114, 114, 112, 115, 111, 111, 112, 117, 117, 113, 115, 111, 193, 193, 189, 199, 130, 195, 196, 195, 201, 196, 198, 189, 148, 114, 114, 121, 122, 156, 152, 147, 145, 132, 133, 140, 174, 156, 107, 106, 115, 125, 122, 157, 164, 159, 153, 144, 128, 129, 128, 123, 109, 111, 111, 122, 128, 150, 137, 113, 128, 155, 155, 135, 157, 147, 179, 187, 191, 193, 193, 192, 198, 195, 197, 197, 199, 193, 192, 182, 176, 154, 150, 146, 159, 168, 192, 192, 197, 201, 203, 205, 208, 206, 205, 200, 192, 192, 162, 161, 143, 155, 138, 163, 218, 230, 231, 231, 231, 230, 230, 230, 231, 231, 229, 228, 230, 231, 231, 231, 227, 228, 228, 229, 228, 229, 224, 226, 224, 227, 228, 222, 228, 224, 228, 226, 225, 223, 223, 222, 222, 224, 224, 222, 222, 222, 222, 220, 220, 208, 162, 143, 139, 141, 130, 132, 132, 130, 131, 131, 132, 128, 117, 117, 117, 116, 115, 112, 112, 107, 112, 119, 118, 114, 115, 117, 108, 109, 108, 108, 113, 111, 105, 123, 122, 107, 107, 109, 109, 113, 105, 106, 106, 108, 108, 130, 120, 117, 116, 114, 116, 116, 132, 122, 117, 118, 128, 123, 121, 129, 118, 122, 112, 118, 111, 110, 109, 112, 112, 107, 103, 107, 110, 124, 125, 131, 112, 116, 118, 126, 124, 119, 122, 120, 118, 115, 122, 121, 117, 123, 121, 124, 124, 123, 122, 126, 122, 131, 125, 124, 119, 124, 117, 116, 117, 116, 122, 120, 113, 115, 119, 112, 124, 115, 115, 116, 116, 114, 197, 191, 191, 193, 112, 186, 194, 199, 193, 195, 194, 188, 148, 111, 112, 121, 129, 165, 162, 160, 153, 132, 136, 149, 168, 162, 113, 109, 129, 128, 114, 148, 165, 160, 152, 141, 134, 134, 137, 131, 115, 108, 113, 110, 113, 135, 137, 115, 136, 157, 155, 140, 160, 149, 178, 193, 193, 191, 189, 196, 193, 196, 193, 198, 197, 194, 194, 189, 180, 165, 156, 150, 158, 166, 187, 192, 193, 198, 198, 204, 206, 206, 206, 196, 194, 195, 165, 168, 146, 153, 144, 166, 223, 228, 229, 230, 231, 229, 229, 230, 227, 231, 230, 230, 229, 229, 231, 231, 226, 227, 228, 230, 231, 228, 222, 226, 223, 223, 224, 225, 224, 222, 224, 225, 225, 222, 222, 223, 221, 224, 226, 221, 221, 225, 216, 224, 219, 210, 166, 141, 140, 134, 132, 135, 132, 130, 133, 130, 135, 125, 127, 122, 118, 113, 118, 116, 116, 117, 117, 124, 119, 120, 120, 123, 121, 111, 118, 120, 117, 117, 115, 116, 118, 113, 112, 109, 110, 112, 114, 113, 109, 108, 108, 129, 120, 121, 124, 123, 126, 124, 133, 124, 124, 118, 124, 126, 128, 134, 120, 118, 118, 110, 116, 110, 113, 110, 112, 111, 108, 112, 109, 126, 122, 133, 115, 117, 122, 124, 122, 123, 121, 124, 121, 121, 125, 120, 118, 126, 127, 132, 125, 122, 128, 125, 131, 126, 124, 128, 122, 129, 117, 119, 121, 124, 121, 130, 124, 127, 117, 122, 125, 122, 128, 126, 122, 115, 192, 190, 194, 192, 113, 186, 195, 193, 194, 194, 197, 184, 146, 122, 112, 128, 132, 162, 167, 164, 157, 138, 145, 163, 182, 169, 121, 129, 127, 127, 116, 146, 148, 155, 142, 137, 132, 128, 140, 138, 121, 115, 110, 117, 122, 130, 138, 120, 143, 157, 155, 141, 155, 149, 177, 190, 196, 195, 189, 193, 195, 190, 193, 199, 196, 195, 192, 190, 177, 169, 158, 159, 157, 163, 187, 194, 197, 197, 202, 202, 202, 202, 198, 192, 192, 186, 171, 166, 144, 152, 152, 165, 222, 228, 231, 230, 231, 229, 229, 229, 230, 230, 229, 230, 229, 229, 230, 228, 226, 229, 227, 228, 230, 226, 222, 223, 224, 226, 226, 227, 224, 225, 224, 226, 225, 225, 220, 222, 224, 226, 225, 226, 221, 224, 222, 220, 219, 210, 172, 148, 142, 145, 140, 133, 137, 135, 138, 131, 133, 135, 129, 129, 118, 115, 116, 120, 122, 116, 120, 122, 122, 125, 117, 115, 118, 116, 123, 122, 120, 115, 116, 125, 123, 120, 112, 117, 119, 115, 117, 117, 116, 119, 115, 126, 131, 128, 124, 120, 125, 119, 122, 124, 126, 118, 128, 124, 121, 137, 127, 121, 114, 112, 114, 112, 112, 112, 117, 107, 107, 114, 113, 124, 131, 134, 123, 124, 127, 128, 134, 129, 126, 122, 123, 125, 128, 127, 122, 125, 129, 130, 127, 126, 132, 128, 130, 128, 125, 131, 126, 132, 126, 123, 128, 130, 130, 127, 126, 125, 122, 123, 128, 123, 122, 123, 116, 120, 194, 187, 190, 196, 109, 187, 191, 195, 191, 191, 193, 186, 142, 123, 111, 124, 132, 161, 168, 170, 162, 162, 167, 178, 183, 172, 145, 132, 126, 133, 121, 137, 138, 140, 131, 124, 118, 116, 137, 128, 121, 124, 116, 121, 122, 123, 143, 124, 143, 161, 153, 142, 152, 148, 178, 193, 194, 192, 197, 193, 193, 199, 192, 199, 198, 193, 195, 189, 177, 170, 156, 156, 157, 166, 178, 190, 197, 197, 200, 202, 203, 203, 200, 193, 192, 188, 167, 156, 142, 162, 147, 168, 219, 227, 231, 231, 231, 230, 230, 229, 229, 230, 229, 228, 229, 230, 230, 226, 226, 225, 219, 225, 229, 227, 226, 222, 224, 224, 224, 224, 222, 223, 223, 221, 223, 222, 220, 223, 222, 221, 224, 222, 219, 219, 221, 217, 219, 211, 184, 149, 147, 143, 146, 143, 145, 145, 140, 138, 140, 135, 142, 134, 128, 128, 121, 127, 122, 124, 124, 126, 132, 128, 122, 123, 117, 122, 129, 123, 121, 116, 122, 125, 126, 126, 121, 118, 119, 123, 122, 119, 119, 124, 123, 127, 132, 133, 127, 127, 128, 122, 134, 121, 121, 119, 125, 129, 127, 142, 124, 128, 116, 118, 116, 117, 129, 117, 115, 117, 112, 111, 121, 124, 135, 129, 119, 128, 128, 129, 135, 131, 127, 134, 125, 129, 128, 126, 127, 132, 130, 129, 132, 127, 126, 132, 129, 129, 128, 131, 135, 131, 130, 127, 123, 129, 130, 126, 126, 125, 126, 123, 125, 122, 121, 124, 116, 118, 193, 187, 189, 193, 116, 191, 192, 193, 195, 194, 184, 184, 145, 119, 110, 127, 143, 167, 169, 169, 169, 173, 172, 180, 181, 177, 146, 131, 126, 136, 123, 132, 133, 134, 124, 116, 120, 119, 132, 135, 123, 130, 123, 123, 125, 124, 140, 126, 147, 158, 154, 142, 155, 151, 177, 190, 196, 192, 194, 192, 192, 199, 198, 200, 197, 194, 191, 188, 170, 168, 158, 157, 159, 164, 173, 190, 192, 198, 199, 202, 201, 200, 198, 190, 188, 184, 165, 155, 150, 159, 155, 168, 224, 229, 231, 231, 230, 229, 230, 228, 228, 229, 228, 230, 229, 228, 228, 227, 225, 225, 228, 225, 228, 227, 226, 221, 224, 224, 223, 223, 225, 223, 223, 223, 223, 222, 221, 220, 222, 222, 222, 216, 220, 216, 216, 221, 216, 210, 185, 158, 154, 151, 151, 150, 150, 152, 150, 142, 150, 141, 147, 140, 132, 132, 123, 127, 129, 127, 122, 126, 128, 129, 127, 124, 119, 118, 125, 126, 128, 121, 119, 131, 132, 129, 132, 123, 124, 121, 129, 127, 137, 135, 125, 130, 138, 130, 120, 130, 125, 131, 138, 134, 126, 126, 137, 133, 129, 149, 134, 131, 121, 121, 123, 123, 124, 120, 116, 119, 114, 118, 119, 130, 134, 130, 121, 129, 128, 131, 133, 131, 128, 131, 132, 135, 135, 131, 136, 128, 134, 134, 133, 133, 135, 136, 134, 133, 130, 133, 136, 132, 128, 128, 131, 132, 128, 129, 128, 127, 122, 126, 120, 125, 126, 125, 126, 122, 186, 188, 188, 192, 111, 188, 192, 197, 193, 192, 190, 182, 139, 111, 111, 128, 144, 169, 168, 171, 166, 172, 177, 182, 187, 183, 147, 120, 133, 120, 115, 121, 125, 126, 121, 119, 114, 119, 127, 135, 118, 127, 122, 131, 122, 125, 144, 129, 143, 155, 150, 145, 154, 154, 178, 192, 195, 196, 190, 194, 194, 196, 195, 195, 197, 196, 198, 191, 179, 173, 160, 157, 158, 161, 167, 178, 195, 196, 199, 198, 198, 202, 192, 190, 191, 176, 160, 155, 148, 160, 155, 170, 221, 228, 228, 228, 229, 228, 229, 230, 229, 229, 228, 229, 229, 228, 229, 226, 226, 227, 229, 226, 227, 228, 225, 224, 224, 224, 224, 223, 226, 220, 226, 223, 221, 220, 219, 220, 221, 221, 221, 223, 222, 219, 216, 221, 216, 214, 195, 162, 163, 162, 157, 156, 156, 153, 155, 157, 150, 147, 149, 143, 130, 131, 128, 128, 133, 129, 128, 126, 126, 131, 131, 130, 123, 120, 131, 127, 132, 135, 131, 135, 128, 128, 130, 128, 135, 132, 128, 123, 136, 130, 132, 127, 135, 136, 126, 133, 134, 136, 134, 137, 131, 128, 136, 142, 130, 142, 137, 137, 129, 130, 131, 134, 131, 127, 126, 118, 121, 124, 125, 132, 141, 142, 128, 130, 138, 140, 137, 134, 135, 138, 136, 133, 137, 137, 133, 135, 138, 135, 138, 130, 134, 137, 133, 131, 135, 141, 136, 134, 135, 134, 130, 136, 124, 130, 127, 129, 124, 127, 125, 121, 122, 128, 129, 124, 190, 190, 188, 193, 116, 193, 195, 194, 189, 188, 189, 179, 135, 113, 122, 122, 146, 165, 163, 170, 168, 172, 180, 184, 185, 186, 149, 130, 134, 114, 120, 116, 125, 118, 119, 117, 125, 119, 130, 135, 124, 125, 127, 126, 129, 126, 144, 133, 141, 166, 159, 146, 156, 155, 184, 189, 197, 191, 194, 189, 192, 193, 192, 197, 196, 195, 194, 194, 183, 171, 165, 159, 160, 164, 168, 168, 196, 199, 196, 199, 199, 197, 191, 190, 190, 179, 159, 157, 151, 160, 155, 177, 218, 226, 229, 228, 227, 227, 226, 228, 229, 229, 226, 226, 228, 230, 229, 227, 226, 225, 227, 228, 227, 224, 222, 222, 223, 222, 227, 225, 224, 224, 224, 228, 223, 219, 220, 220, 223, 222, 221, 220, 221, 218, 216, 221, 218, 208, 202, 173, 170, 168, 165, 161, 158, 155, 152, 154, 152, 149, 153, 146, 140, 138, 131, 137, 133, 127, 132, 129, 132, 127, 128, 131, 125, 124, 132, 128, 125, 135, 134, 135, 129, 134, 134, 131, 133, 130, 128, 126, 130, 128, 128, 135, 136, 136, 128, 134, 132, 139, 143, 130, 134, 136, 140, 149, 140, 147, 143, 139, 136, 135, 147, 144, 131, 130, 125, 131, 129, 127, 135, 130, 140, 142, 135, 136, 136, 133, 137, 137, 132, 135, 134, 136, 134, 138, 133, 140, 141, 140, 138, 144, 144, 141, 140, 138, 137, 141, 141, 129, 132, 131, 129, 133, 134, 132, 134, 133, 130, 135, 129, 135, 122, 134, 127, 131, 189, 190, 187, 186, 119, 186, 191, 190, 189, 191, 185, 179, 133, 120, 119, 128, 144, 162, 169, 168, 171, 173, 186, 185, 192, 187, 144, 135, 122, 115, 119, 121, 122, 119, 125, 127, 127, 124, 135, 130, 126, 132, 131, 127, 132, 133, 142, 136, 147, 169, 167, 148, 160, 159, 187, 191, 196, 194, 196, 191, 197, 198, 199, 199, 199, 193, 192, 196, 186, 176, 166, 157, 162, 164, 168, 170, 193, 198, 195, 197, 197, 187, 182, 189, 189, 179, 157, 160, 153, 158, 156, 169, 218, 224, 226, 228, 228, 227, 224, 225, 227, 228, 227, 226, 227, 229, 227, 227, 224, 223, 224, 225, 226, 224, 222, 223, 224, 225, 224, 221, 221, 223, 220, 224, 217, 217, 221, 221, 223, 221, 222, 215, 215, 218, 221, 216, 215, 208, 196, 176, 183, 184, 183, 169, 171, 166, 161, 156, 159, 154, 155, 147, 148, 139, 138, 138, 135, 134, 136, 135, 137, 133, 134, 128, 126, 129, 133, 133, 134, 135, 130, 136, 137, 135, 129, 137, 133, 135, 139, 137, 136, 134, 139, 139, 142, 140, 140, 142, 145, 136, 145, 133, 134, 140, 146, 147, 137, 144, 143, 143, 139, 136, 133, 131, 126, 134, 132, 129, 129, 129, 132, 133, 144, 139, 132, 134, 140, 136, 140, 133, 139, 136, 139, 136, 137, 141, 139, 145, 144, 141, 139, 147, 145, 146, 140, 137, 142, 139, 143, 137, 139, 135, 138, 139, 133, 134, 135, 130, 133, 133, 131, 131, 129, 132, 128, 128, 188, 187, 186, 187, 95, 183, 191, 191, 190, 191, 191, 183, 131, 125, 121, 126, 145, 163, 165, 169, 170, 175, 181, 185, 187, 181, 163, 138, 122, 119, 121, 121, 123, 128, 124, 128, 139, 128, 139, 137, 134, 125, 135, 134, 138, 136, 143, 133, 145, 171, 167, 151, 162, 154, 186, 193, 190, 194, 192, 192, 194, 192, 193, 193, 194, 196, 191, 190, 181, 176, 170, 166, 164, 168, 169, 172, 195, 197, 197, 195, 196, 185, 181, 180, 186, 172, 161, 159, 153, 162, 156, 169, 218, 225, 228, 228, 227, 225, 225, 226, 227, 225, 226, 226, 226, 229, 226, 226, 221, 223, 224, 225, 225, 221, 220, 221, 223, 224, 224, 222, 222, 220, 221, 223, 219, 219, 217, 218, 222, 221, 218, 217, 217, 219, 216, 214, 214, 209, 200, 195, 203, 207, 196, 190, 193, 184, 182, 173, 168, 164, 164, 156, 155, 146, 143, 140, 143, 139, 138, 142, 136, 141, 146, 135, 134, 138, 139, 142, 139, 136, 137, 138, 136, 141, 129, 129, 128, 137, 139, 142, 144, 142, 140, 142, 143, 143, 145, 143, 151, 151, 149, 142, 140, 140, 140, 148, 137, 143, 144, 143, 137, 139, 129, 134, 128, 133, 132, 134, 130, 134, 131, 141, 145, 136, 134, 141, 141, 144, 136, 139, 138, 135, 139, 137, 143, 142, 140, 143, 143, 143, 146, 140, 141, 144, 137, 136, 143, 140, 140, 142, 144, 141, 142, 144, 136, 144, 143, 138, 136, 136, 143, 131, 135, 132, 130, 133, 189, 186, 185, 183, 91, 177, 195, 192, 191, 190, 186, 179, 133, 123, 114, 121, 142, 153, 159, 163, 166, 173, 182, 183, 186, 181, 174, 134, 122, 119, 124, 125, 122, 125, 129, 135, 130, 130, 136, 138, 135, 136, 138, 136, 135, 131, 144, 138, 145, 169, 164, 153, 162, 158, 182, 190, 194, 195, 194, 189, 194, 194, 195, 199, 198, 197, 191, 193, 178, 175, 176, 163, 170, 174, 170, 177, 196, 198, 196, 195, 189, 184, 171, 171, 172, 168, 161, 158, 155, 163, 152, 174, 213, 224, 226, 227, 226, 227, 228, 226, 226, 224, 225, 224, 227, 227, 229, 228, 224, 223, 222, 224, 222, 220, 217, 217, 221, 221, 222, 223, 221, 220, 219, 219, 218, 218, 211, 214, 219, 220, 216, 215, 214, 218, 219, 213, 215, 215, 212, 209, 207, 203, 201, 201, 204, 201, 197, 198, 193, 192, 184, 175, 170, 164, 160, 151, 141, 146, 143, 145, 146, 144, 144, 145, 139, 141, 139, 144, 142, 136, 138, 139, 140, 147, 139, 134, 135, 140, 137, 137, 137, 140, 138, 143, 147, 145, 140, 144, 153, 151, 146, 147, 145, 144, 148, 153, 143, 144, 142, 148, 135, 138, 137, 136, 139, 135, 140, 132, 134, 134, 134, 135, 144, 144, 139, 140, 147, 138, 143, 140, 142, 142, 144, 143, 147, 147, 143, 143, 143, 142, 146, 141, 142, 148, 138, 145, 149, 143, 143, 146, 147, 140, 140, 141, 141, 144, 144, 142, 136, 139, 144, 141, 135, 138, 135, 135, 186, 182, 181, 183, 91, 178, 184, 188, 189, 192, 182, 177, 141, 128, 124, 132, 142, 159, 142, 147, 153, 164, 179, 184, 183, 179, 172, 130, 123, 119, 126, 127, 129, 133, 130, 131, 134, 128, 137, 137, 138, 144, 139, 136, 131, 133, 144, 140, 145, 171, 169, 160, 169, 157, 181, 188, 188, 193, 190, 194, 192, 194, 191, 198, 194, 188, 193, 193, 184, 176, 176, 174, 171, 176, 173, 192, 196, 195, 193, 192, 188, 177, 166, 168, 169, 166, 163, 160, 157, 167, 156, 176, 215, 214, 223, 226, 226, 226, 227, 226, 227, 224, 222, 226, 227, 228, 226, 225, 224, 223, 223, 222, 223, 218, 216, 220, 220, 222, 221, 220, 219, 219, 220, 221, 218, 214, 213, 215, 215, 217, 214, 217, 217, 219, 217, 215, 215, 216, 211, 209, 211, 204, 205, 201, 206, 204, 202, 202, 200, 202, 199, 198, 195, 185, 182, 174, 159, 148, 145, 144, 146, 143, 146, 143, 146, 142, 143, 147, 145, 141, 141, 145, 140, 146, 137, 135, 137, 139, 142, 143, 141, 146, 143, 138, 147, 141, 144, 144, 154, 156, 147, 152, 151, 146, 150, 153, 148, 146, 147, 149, 143, 141, 141, 142, 139, 140, 144, 142, 139, 139, 139, 138, 143, 141, 144, 140, 142, 146, 149, 146, 141, 151, 149, 152, 145, 147, 143, 148, 145, 148, 143, 145, 148, 145, 147, 138, 148, 136, 148, 143, 146, 141, 140, 143, 142, 141, 140, 142, 141, 138, 139, 144, 136, 141, 136, 134, 184, 187, 183, 188, 97, 174, 185, 186, 186, 189, 184, 173, 141, 127, 120, 134, 139, 148, 140, 142, 145, 154, 175, 182, 185, 181, 172, 128, 125, 126, 130, 127, 134, 131, 133, 133, 133, 135, 136, 142, 136, 140, 138, 138, 136, 138, 145, 141, 148, 171, 158, 160, 164, 158, 182, 188, 189, 195, 193, 188, 197, 193, 191, 197, 194, 193, 197, 193, 186, 178, 177, 177, 170, 180, 180, 195, 192, 192, 193, 189, 182, 180, 166, 166, 172, 169, 164, 160, 158, 163, 165, 178, 213, 217, 221, 226, 227, 222, 224, 226, 226, 225, 225, 223, 225, 226, 223, 223, 223, 222, 222, 222, 224, 221, 218, 220, 220, 220, 220, 221, 218, 220, 220, 221, 219, 220, 214, 217, 214, 215, 217, 216, 215, 219, 216, 217, 211, 215, 212, 212, 214, 207, 207, 203, 202, 204, 201, 205, 203, 203, 202, 203, 195, 193, 192, 184, 172, 163, 156, 155, 144, 151, 150, 151, 149, 147, 147, 149, 144, 145, 143, 143, 145, 144, 138, 141, 144, 147, 146, 151, 143, 146, 147, 149, 152, 151, 145, 150, 160, 154, 154, 152, 154, 148, 151, 147, 148, 146, 150, 152, 149, 145, 145, 141, 142, 148, 143, 143, 140, 144, 145, 144, 145, 142, 142, 145, 147, 151, 150, 148, 149, 151, 151, 152, 147, 152, 148, 152, 149, 149, 155, 147, 148, 149, 152, 146, 150, 145, 146, 144, 152, 148, 147, 149, 147, 149, 147, 143, 143, 141, 147, 147, 143, 145, 144, 140, 186, 184, 183, 192, 97, 180, 185, 187, 189, 187, 187, 170, 140, 130, 123, 128, 140, 149, 145, 147, 142, 150, 169, 180, 179, 176, 170, 143, 129, 134, 129, 131, 135, 129, 131, 133, 129, 131, 143, 140, 141, 143, 146, 136, 140, 138, 144, 143, 153, 169, 160, 157, 158, 161, 180, 187, 190, 190, 194, 193, 196, 195, 195, 194, 197, 195, 192, 192, 188, 182, 178, 180, 172, 177, 183, 191, 193, 198, 195, 187, 181, 174, 169, 171, 172, 168, 166, 163, 163, 165, 163, 178, 210, 221, 218, 223, 225, 225, 225, 226, 227, 228, 225, 226, 225, 224, 224, 223, 222, 220, 223, 219, 220, 222, 219, 221, 220, 222, 220, 221, 218, 218, 219, 220, 220, 219, 216, 217, 218, 217, 215, 216, 216, 216, 217, 214, 213, 214, 211, 214, 209, 209, 205, 208, 200, 205, 206, 206, 204, 203, 200, 201, 198, 198, 189, 179, 170, 165, 162, 154, 155, 156, 154, 159, 159, 149, 159, 151, 154, 150, 147, 144, 150, 149, 147, 145, 144, 147, 151, 148, 145, 147, 147, 147, 149, 148, 143, 153, 148, 146, 150, 150, 148, 146, 148, 151, 151, 148, 151, 148, 150, 143, 144, 144, 140, 150, 147, 144, 145, 147, 143, 150, 151, 146, 147, 147, 146, 151, 156, 152, 146, 144, 152, 153, 148, 155, 152, 152, 152, 154, 150, 151, 153, 152, 157, 155, 153, 150, 154, 151, 154, 151, 150, 154, 151, 155, 153, 146, 149, 148, 147, 146, 148, 155, 152, 146, 186, 181, 184, 184, 93, 173, 186, 187, 188, 188, 184, 175, 143, 134, 128, 130, 142, 149, 150, 151, 144, 151, 165, 172, 174, 173, 170, 141, 127, 136, 137, 134, 135, 136, 134, 135, 139, 140, 150, 145, 147, 144, 144, 141, 137, 144, 148, 142, 146, 167, 163, 156, 165, 165, 182, 185, 193, 195, 194, 197, 194, 194, 196, 194, 196, 198, 192, 199, 184, 182, 170, 170, 168, 172, 175, 183, 190, 193, 186, 181, 177, 171, 166, 166, 175, 168, 168, 164, 160, 175, 165, 183, 208, 220, 219, 225, 223, 226, 227, 225, 227, 229, 227, 226, 223, 225, 224, 223, 223, 222, 220, 218, 222, 219, 220, 220, 224, 222, 221, 224, 218, 217, 217, 219, 218, 218, 218, 218, 219, 219, 216, 217, 221, 218, 220, 215, 213, 214, 212, 214, 209, 212, 208, 208, 208, 207, 209, 204, 211, 202, 203, 200, 196, 193, 180, 168, 170, 164, 161, 161, 161, 162, 163, 163, 167, 152, 156, 156, 155, 149, 153, 149, 153, 152, 149, 148, 149, 155, 156, 153, 154, 149, 147, 150, 150, 153, 149, 157, 154, 152, 153, 149, 152, 149, 151, 152, 150, 143, 152, 149, 151, 147, 151, 147, 147, 150, 149, 151, 150, 147, 149, 152, 149, 148, 153, 146, 153, 154, 156, 147, 153, 155, 151, 152, 154, 149, 149, 153, 155, 158, 156, 154, 155, 153, 155, 153, 151, 154, 151, 155, 153, 154, 154, 155, 154, 158, 157, 154, 154, 154, 150, 151, 150, 156, 152, 147, 186, 185, 182, 185, 87, 180, 190, 190, 190, 187, 181, 177, 139, 131, 128, 131, 140, 145, 142, 147, 142, 149, 148, 168, 171, 168, 167, 149, 131, 132, 136, 132, 137, 142, 138, 142, 145, 142, 154, 150, 152, 150, 145, 145, 143, 144, 152, 147, 153, 171, 163, 161, 169, 169, 185, 190, 196, 195, 194, 196, 195, 198, 197, 195, 196, 202, 195, 196, 188, 179, 169, 161, 165, 167, 170, 177, 184, 184, 181, 180, 173, 171, 166, 169, 172, 167, 164, 165, 166, 175, 166, 181, 211, 221, 221, 225, 224, 223, 225, 225, 226, 226, 226, 227, 222, 225, 224, 222, 220, 222, 221, 220, 223, 221, 219, 219, 221, 221, 221, 220, 219, 219, 219, 221, 217, 218, 214, 219, 219, 221, 215, 219, 217, 217, 221, 218, 214, 216, 216, 214, 212, 210, 209, 207, 206, 212, 210, 208, 209, 200, 198, 198, 192, 180, 176, 169, 170, 162, 161, 159, 162, 167, 164, 169, 163, 159, 156, 162, 152, 156, 156, 155, 162, 158, 156, 157, 148, 156, 155, 158, 152, 151, 156, 155, 151, 161, 156, 154, 153, 156, 155, 152, 146, 149, 145, 157, 157, 149, 153, 152, 158, 150, 151, 148, 153, 152, 152, 151, 150, 149, 149, 151, 155, 151, 156, 143, 155, 155, 153, 153, 152, 158, 153, 151, 155, 150, 154, 154, 149, 154, 155, 159, 157, 163, 158, 157, 156, 157, 158, 155, 156, 152, 154, 155, 159, 161, 159, 157, 158, 157, 155, 155, 162, 168, 161, 156, 188, 182, 184, 187, 88, 178, 192, 189, 190, 192, 181, 170, 142, 130, 132, 130, 130, 140, 137, 139, 144, 138, 148, 157, 161, 159, 154, 147, 141, 138, 139, 138, 136, 136, 140, 145, 144, 143, 151, 149, 154, 149, 148, 150, 146, 147, 152, 149, 157, 173, 168, 166, 171, 174, 186, 192, 195, 192, 192, 193, 197, 199, 196, 200, 196, 204, 197, 195, 186, 171, 168, 165, 171, 166, 166, 173, 177, 180, 177, 181, 174, 173, 170, 173, 170, 172, 173, 169, 170, 170, 168, 181, 213, 224, 222, 224, 225, 225, 222, 224, 226, 223, 228, 224, 225, 225, 222, 222, 220, 218, 223, 223, 223, 221, 220, 222, 222, 223, 224, 221, 218, 220, 221, 221, 218, 219, 218, 218, 222, 220, 219, 219, 218, 216, 216, 217, 216, 215, 214, 214, 208, 208, 213, 208, 210, 213, 210, 205, 205, 201, 197, 190, 185, 177, 178, 172, 170, 167, 167, 165, 168, 171, 170, 173, 168, 167, 161, 165, 160, 162, 159, 165, 162, 165, 158, 155, 151, 156, 160, 154, 153, 153, 157, 159, 158, 157, 156, 160, 153, 163, 153, 157, 152, 153, 151, 155, 157, 153, 155, 158, 155, 154, 151, 152, 149, 153, 151, 153, 154, 156, 151, 152, 153, 157, 154, 150, 149, 159, 159, 156, 156, 158, 158, 159, 156, 157, 153, 156, 158, 161, 158, 160, 162, 163, 162, 165, 161, 159, 165, 164, 162, 160, 158, 163, 158, 159, 160, 161, 157, 166, 155, 163, 165, 168, 163, 161, 184, 185, 182, 184, 87, 182, 190, 187, 191, 190, 181, 170, 142, 133, 132, 130, 134, 138, 140, 140, 137, 138, 150, 151, 154, 153, 144, 145, 140, 136, 136, 142, 134, 137, 137, 142, 147, 147, 149, 157, 149, 147, 147, 146, 153, 151, 151, 157, 156, 173, 170, 164, 172, 175, 190, 195, 199, 193, 194, 192, 198, 196, 195, 198, 196, 199, 195, 197, 190, 177, 171, 169, 171, 171, 170, 170, 172, 176, 181, 176, 173, 174, 174, 176, 173, 174, 171, 169, 173, 178, 169, 186, 214, 221, 222, 226, 221, 223, 225, 225, 225, 226, 226, 225, 224, 224, 224, 221, 220, 220, 220, 221, 222, 219, 222, 221, 222, 223, 224, 219, 219, 219, 220, 218, 220, 218, 216, 220, 221, 218, 219, 218, 219, 217, 216, 219, 217, 215, 215, 211, 214, 211, 211, 208, 210, 211, 211, 209, 207, 203, 198, 188, 178, 177, 172, 169, 172, 171, 172, 170, 174, 178, 179, 171, 175, 169, 170, 164, 164, 163, 163, 160, 163, 161, 163, 161, 159, 163, 163, 158, 163, 156, 159, 161, 160, 157, 157, 157, 159, 154, 159, 155, 155, 158, 163, 156, 158, 157, 157, 160, 156, 158, 155, 156, 157, 154, 156, 154, 158, 152, 154, 152, 158, 156, 151, 156, 154, 155, 157, 157, 160, 160, 160, 159, 160, 158, 162, 154, 162, 162, 162, 162, 167, 167, 162, 169, 166, 161, 167, 168, 165, 164, 160, 159, 162, 161, 161, 159, 164, 160, 161, 164, 165, 166, 159, 157, 189, 182, 179, 181, 80, 181, 189, 191, 190, 190, 180, 169, 147, 138, 136, 136, 139, 139, 143, 139, 140, 145, 151, 157, 156, 159, 151, 155, 140, 141, 131, 138, 134, 140, 141, 146, 147, 146, 147, 150, 153, 146, 147, 154, 146, 153, 153, 155, 162, 178, 172, 172, 176, 179, 193, 194, 200, 197, 199, 193, 195, 193, 193, 199, 199, 194, 197, 195, 188, 177, 177, 170, 178, 174, 175, 173, 172, 181, 180, 179, 172, 176, 173, 174, 177, 170, 169, 173, 168, 176, 172, 185, 212, 221, 220, 225, 220, 226, 226, 225, 225, 225, 223, 223, 220, 223, 220, 222, 221, 221, 220, 221, 221, 221, 220, 222, 222, 221, 223, 219, 219, 217, 219, 219, 217, 217, 216, 216, 217, 219, 216, 215, 215, 216, 213, 217, 215, 212, 216, 211, 212, 208, 211, 209, 213, 213, 210, 209, 204, 196, 194, 188, 180, 180, 179, 178, 176, 174, 178, 178, 174, 176, 178, 173, 174, 167, 175, 168, 165, 165, 166, 170, 167, 167, 164, 159, 165, 163, 161, 161, 164, 161, 159, 160, 160, 158, 159, 161, 159, 158, 163, 163, 163, 160, 164, 161, 161, 160, 159, 161, 154, 158, 150, 157, 157, 157, 157, 159, 152, 155, 153, 152, 156, 159, 158, 157, 153, 160, 162, 157, 157, 160, 159, 161, 161, 160, 161, 166, 163, 166, 169, 168, 172, 168, 167, 168, 167, 166, 167, 174, 171, 166, 165, 164, 164, 164, 162, 162, 167, 168, 170, 165, 168, 164, 169, 157, 187, 182, 176, 179, 78, 181, 182, 186, 186, 190, 185, 167, 145, 141, 141, 139, 138, 144, 147, 145, 148, 148, 163, 166, 166, 163, 159, 155, 146, 139, 134, 138, 140, 144, 145, 150, 149, 146, 148, 155, 155, 153, 155, 151, 153, 153, 154, 151, 162, 172, 167, 175, 175, 176, 192, 196, 198, 198, 194, 198, 193, 197, 199, 198, 195, 198, 196, 195, 187, 175, 178, 172, 174, 177, 172, 169, 169, 172, 182, 176, 168, 169, 172, 174, 174, 170, 171, 172, 172, 177, 177, 190, 211, 220, 220, 222, 220, 225, 225, 224, 225, 224, 225, 221, 220, 224, 222, 220, 218, 219, 219, 219, 223, 221, 219, 220, 219, 220, 220, 218, 214, 216, 215, 217, 219, 219, 218, 218, 218, 218, 216, 214, 216, 214, 213, 214, 215, 214, 212, 214, 214, 213, 213, 212, 213, 213, 209, 208, 202, 195, 191, 186, 185, 178, 174, 176, 177, 178, 179, 184, 180, 177, 183, 177, 178, 170, 175, 176, 172, 163, 169, 166, 166, 172, 162, 163, 161, 161, 168, 169, 168, 165, 159, 159, 163, 163, 161, 160, 161, 161, 163, 164, 162, 160, 159, 159, 162, 160, 161, 166, 161, 158, 158, 154, 160, 163, 165, 159, 153, 159, 155, 152, 163, 161, 159, 157, 160, 164, 163, 166, 162, 161, 165, 164, 160, 161, 161, 167, 164, 164, 166, 166, 172, 173, 173, 168, 168, 168, 168, 171, 165, 168, 166, 169, 165, 164, 162, 164, 166, 168, 166, 167, 168, 169, 171, 162, 184, 184, 183, 182, 81, 182, 190, 188, 187, 188, 182, 163, 140, 145, 144, 141, 146, 153, 157, 154, 154, 159, 161, 174, 170, 167, 163, 149, 151, 143, 138, 144, 138, 142, 144, 150, 153, 151, 153, 156, 162, 158, 151, 150, 153, 155, 156, 157, 161, 177, 170, 173, 181, 178, 194, 199, 193, 196, 191, 195, 189, 197, 200, 201, 199, 199, 195, 198, 184, 174, 177, 171, 174, 171, 171, 171, 170, 171, 178, 180, 171, 174, 172, 178, 179, 178, 176, 179, 180, 179, 181, 193, 211, 216, 217, 221, 218, 221, 224, 223, 226, 225, 225, 222, 219, 220, 214, 219, 219, 218, 218, 217, 220, 220, 220, 220, 219, 223, 221, 217, 216, 215, 215, 216, 217, 216, 214, 220, 217, 219, 215, 214, 216, 217, 213, 215, 216, 216, 211, 213, 212, 212, 214, 206, 215, 212, 206, 206, 201, 197, 187, 183, 180, 181, 178, 182, 181, 181, 181, 183, 180, 184, 179, 177, 178, 172, 175, 179, 176, 166, 163, 167, 167, 165, 172, 166, 168, 169, 170, 171, 163, 165, 162, 164, 166, 163, 157, 161, 163, 165, 163, 163, 162, 163, 162, 167, 167, 164, 166, 158, 165, 157, 159, 162, 158, 163, 160, 162, 157, 163, 159, 160, 158, 158, 157, 163, 161, 161, 160, 162, 158, 165, 161, 163, 158, 160, 162, 164, 163, 164, 165, 166, 171, 172, 171, 164, 170, 167, 168, 172, 168, 170, 164, 167, 165, 160, 167, 158, 163, 164, 168, 170, 173, 172, 166, 159, 189, 183, 176, 180, 74, 177, 186, 186, 188, 187, 183, 164, 145, 148, 141, 144, 149, 154, 156, 158, 162, 160, 172, 172, 170, 169, 154, 146, 150, 148, 142, 143, 143, 149, 149, 147, 151, 146, 157, 157, 160, 155, 156, 155, 157, 158, 159, 159, 167, 176, 172, 173, 181, 179, 189, 196, 191, 198, 193, 194, 195, 193, 198, 197, 198, 201, 198, 195, 190, 174, 178, 179, 174, 174, 166, 169, 175, 168, 181, 176, 174, 182, 182, 174, 181, 181, 174, 179, 179, 178, 180, 192, 215, 216, 220, 221, 222, 220, 222, 224, 225, 224, 223, 222, 221, 220, 218, 219, 218, 217, 218, 218, 220, 222, 219, 221, 220, 222, 217, 214, 214, 216, 215, 218, 217, 219, 217, 220, 218, 217, 214, 215, 216, 216, 217, 214, 213, 214, 214, 213, 215, 216, 213, 214, 214, 211, 210, 206, 202, 192, 187, 184, 185, 182, 181, 183, 181, 184, 185, 183, 185, 183, 183, 182, 177, 174, 182, 179, 182, 170, 170, 168, 172, 174, 176, 171, 173, 175, 169, 175, 165, 168, 165, 167, 169, 164, 163, 168, 165, 164, 170, 165, 169, 170, 175, 173, 171, 168, 171, 162, 169, 163, 167, 169, 161, 161, 161, 162, 162, 158, 162, 158, 161, 162, 162, 161, 163, 156, 165, 158, 157, 164, 159, 162, 155, 156, 160, 160, 165, 160, 163, 165, 166, 172, 172, 167, 171, 168, 172, 168, 171, 167, 164, 170, 169, 170, 160, 168, 169, 172, 169, 176, 171, 170, 170, 161, 185, 182, 177, 185, 80, 184, 188, 190, 188, 186, 184, 160, 150, 148, 144, 150, 153, 157, 163, 161, 164, 161, 175, 171, 167, 172, 156, 153, 159, 149, 146, 144, 149, 151, 152, 151, 150, 153, 154, 162, 159, 161, 162, 161, 165, 157, 162, 163, 163, 176, 171, 173, 179, 179, 188, 193, 194, 190, 191, 193, 191, 190, 197, 198, 198, 198, 195, 194, 188, 179, 178, 179, 176, 172, 173, 174, 176, 173, 180, 179, 179, 180, 181, 183, 182, 184, 172, 180, 179, 179, 179, 188, 212, 216, 219, 217, 222, 219, 223, 222, 224, 221, 222, 218, 222, 221, 220, 220, 217, 216, 216, 218, 222, 221, 216, 217, 220, 219, 220, 218, 214, 218, 217, 219, 217, 218, 214, 214, 216, 218, 215, 215, 217, 215, 215, 211, 216, 214, 216, 213, 212, 215, 216, 209, 211, 209, 206, 203, 201, 190, 186, 187, 181, 183, 184, 180, 180, 182, 185, 183, 183, 181, 180, 181, 177, 177, 180, 173, 179, 182, 170, 172, 171, 174, 180, 177, 171, 172, 175, 167, 169, 172, 166, 169, 170, 168, 170, 170, 170, 175, 172, 173, 175, 176, 176, 174, 177, 175, 173, 175, 172, 175, 171, 168, 166, 167, 165, 165, 161, 157, 158, 160, 163, 159, 162, 162, 165, 163, 164, 162, 157, 155, 161, 156, 150, 159, 161, 163, 165, 164, 166, 172, 173, 174, 174, 170, 170, 168, 172, 172, 180, 177, 177, 181, 176, 178, 176, 180, 180, 184, 181, 181, 178, 179, 179, 175, 178, 180, 180, 184, 89, 181, 189, 184, 188, 187, 182, 161, 150, 144, 145, 150, 154, 160, 167, 165, 167, 168, 171, 170, 171, 162, 157, 154, 157, 154, 150, 150, 147, 152, 148, 154, 155, 156, 162, 166, 166, 167, 168, 174, 173, 168, 163, 165, 167, 177, 176, 174, 183, 181, 185, 191, 193, 192, 186, 192, 189, 188, 193, 199, 196, 195, 196, 193, 189, 178, 176, 173, 174, 168, 175, 170, 176, 174, 177, 177, 186, 182, 188, 180, 185, 181, 179, 181, 183, 185, 178, 192, 210, 213, 220, 221, 222, 220, 221, 220, 223, 221, 220, 221, 220, 220, 220, 216, 215, 216, 220, 221, 220, 218, 212, 216, 215, 215, 219, 215, 216, 214, 218, 218, 215, 213, 216, 214, 212, 218, 214, 215, 213, 215, 215, 216, 215, 213, 213, 216, 214, 209, 211, 210, 210, 210, 206, 202, 190, 189, 191, 188, 188, 186, 182, 183, 181, 185, 184, 181, 186, 185, 180, 180, 180, 173, 176, 174, 176, 181, 177, 167, 171, 177, 170, 176, 172, 173, 171, 171, 168, 173, 170, 176, 174, 171, 171, 172, 179, 177, 177, 174, 179, 176, 182, 180, 176, 177, 173, 175, 174, 171, 170, 171, 166, 170, 163, 165, 158, 157, 163, 164, 162, 160, 162, 164, 167, 163, 162, 164, 162, 162, 165, 162, 157, 163, 164, 166, 174, 178, 177, 179, 180, 181, 180, 181, 184, 182, 183, 186, 189, 185, 187, 187, 185, 185, 190, 187, 190, 190, 187, 187, 187, 188, 185, 179, 182, 178, 174, 182, 71, 180, 185, 187, 184, 183, 177, 160, 151, 150, 150, 153, 160, 166, 164, 165, 169, 168, 172, 170, 167, 168, 153, 155, 153, 155, 152, 149, 152, 152, 154, 153, 168, 166, 166, 175, 177, 177, 177, 178, 179, 171, 166, 165, 169, 175, 173, 175, 182, 183, 191, 188, 192, 186, 186, 186, 189, 190, 194, 198, 192, 195, 193, 197, 190, 175, 178, 174, 176, 169, 173, 172, 174, 179, 180, 183, 183, 182, 187, 180, 179, 185, 175, 180, 181, 186, 183, 194, 209, 212, 218, 221, 220, 218, 220, 222, 221, 220, 221, 217, 218, 217, 219, 218, 213, 216, 218, 221, 216, 215, 216, 212, 213, 213, 213, 210, 213, 214, 217, 218, 215, 214, 217, 215, 214, 215, 214, 208, 214, 219, 214, 215, 215, 214, 212, 213, 216, 211, 208, 211, 211, 206, 205, 194, 187, 183, 189, 188, 188, 187, 184, 185, 181, 187, 184, 184, 186, 181, 184, 184, 182, 176, 177, 176, 177, 175, 174, 171, 176, 172, 172, 171, 172, 173, 175, 172, 171, 173, 175, 176, 176, 179, 177, 178, 175, 176, 176, 173, 173, 173, 177, 175, 176, 176, 172, 174, 170, 169, 168, 171, 168, 171, 170, 170, 167, 162, 165, 167, 168, 160, 160, 164, 167, 167, 165, 161, 164, 163, 164, 164, 168, 169, 172, 184, 184, 188, 192, 193, 189, 193, 193, 192, 194, 189, 186, 194, 199, 190, 195, 199, 201, 202, 202, 205, 206, 204, 205, 203, 206, 207, 206, 207, 197, 192, 189, 202, 115, 192, 188, 185, 178, 175, 180, 166, 158, 156, 160, 154, 159, 166, 167, 166, 161, 166, 170, 168, 171, 165, 154, 158, 162, 158, 150, 149, 151, 151, 153, 157, 162, 161, 165, 166, 174, 169, 167, 172, 173, 169, 161, 163, 169, 170, 169, 174, 176, 172, 180, 181, 179, 181, 180, 171, 178, 179, 183, 186, 186, 185, 188, 184, 177, 166, 166, 154, 161, 163, 158, 162, 165, 163, 169, 170, 169, 168, 172, 169, 171, 172, 163, 163, 169, 173, 175, 181, 194, 192, 192, 200, 198, 195, 202, 200, 201, 202, 200, 198, 200, 201, 196, 197, 194, 195, 198, 197, 207, 202, 198, 201, 193, 189, 191, 183, 190, 189, 190, 192, 192, 192, 192, 188, 187, 185, 187, 186, 196, 206, 199, 194, 193, 188, 192, 190, 192, 194, 193, 199, 203, 210, 213, 211, 206, 190, 208, 191, 190, 185, 192, 199, 195, 179, 180, 177, 174, 164, 188, 177, 172, 159, 152, 152, 148, 153, 144, 148, 156, 160, 172, 160, 157, 160, 164, 163, 170, 161, 161, 193, 187, 196, 189, 204, 206, 187, 176, 193, 170, 154, 139, 138, 139, 140, 135, 158, 149, 149, 147, 160, 142, 153, 166, 140, 147, 150, 137, 154, 166, 148, 133, 131, 133, 134, 152, 136, 137, 151, 139, 134, 136, 137, 132, 141, 145, 146, 150, 151, 147, 149, 149, 159, 156, 163, 188, 163, 151, 144, 141, 140, 155, 134, 130, 146, 131, 152, 147, 140, 137, 142, 155, 159);

begin
process (clk) 
begin
if clk'event and clk = '1' then
 if cs = '1' then
 -- if we = '1' then
  -- memory(address)<= data_in;--memory(to_integer(unsigned(address))) <= data_in;
  -- data_out <= data_in;
  --else
  data_out <= memory(address);
--data_out <= memory(to_integer(unsigned(address)));
  --end if;
 end if;
end if;
end process;
end Behavioral;